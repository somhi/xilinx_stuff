
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"38",x"78",x"00",x"42"),
     1 => (x"6c",x"c6",x"c2",x"6a"),
     2 => (x"00",x"60",x"00",x"38"),
     3 => (x"00",x"00",x"60",x"00"),
     4 => (x"5e",x"0e",x"00",x"60"),
     5 => (x"0e",x"5d",x"5c",x"5b"),
     6 => (x"c2",x"4c",x"71",x"1e"),
     7 => (x"4d",x"bf",x"f2",x"ef"),
     8 => (x"1e",x"c0",x"4b",x"c0"),
     9 => (x"c7",x"02",x"ab",x"74"),
    10 => (x"48",x"a6",x"c4",x"87"),
    11 => (x"87",x"c5",x"78",x"c0"),
    12 => (x"c1",x"48",x"a6",x"c4"),
    13 => (x"1e",x"66",x"c4",x"78"),
    14 => (x"df",x"ee",x"49",x"73"),
    15 => (x"c0",x"86",x"c8",x"87"),
    16 => (x"ef",x"ef",x"49",x"e0"),
    17 => (x"4a",x"a5",x"c4",x"87"),
    18 => (x"f0",x"f0",x"49",x"6a"),
    19 => (x"87",x"c6",x"f1",x"87"),
    20 => (x"83",x"c1",x"85",x"cb"),
    21 => (x"04",x"ab",x"b7",x"c8"),
    22 => (x"26",x"87",x"c7",x"ff"),
    23 => (x"4c",x"26",x"4d",x"26"),
    24 => (x"4f",x"26",x"4b",x"26"),
    25 => (x"c2",x"4a",x"71",x"1e"),
    26 => (x"c2",x"5a",x"f6",x"ef"),
    27 => (x"c7",x"48",x"f6",x"ef"),
    28 => (x"dd",x"fe",x"49",x"78"),
    29 => (x"1e",x"4f",x"26",x"87"),
    30 => (x"4a",x"71",x"1e",x"73"),
    31 => (x"03",x"aa",x"b7",x"c0"),
    32 => (x"cf",x"c2",x"87",x"d3"),
    33 => (x"c4",x"05",x"bf",x"fe"),
    34 => (x"c2",x"4b",x"c1",x"87"),
    35 => (x"c2",x"4b",x"c0",x"87"),
    36 => (x"c4",x"5b",x"c2",x"d0"),
    37 => (x"c2",x"d0",x"c2",x"87"),
    38 => (x"fe",x"cf",x"c2",x"5a"),
    39 => (x"9a",x"c1",x"4a",x"bf"),
    40 => (x"49",x"a2",x"c0",x"c1"),
    41 => (x"fc",x"87",x"e8",x"ec"),
    42 => (x"fe",x"cf",x"c2",x"48"),
    43 => (x"ef",x"fe",x"78",x"bf"),
    44 => (x"4a",x"71",x"1e",x"87"),
    45 => (x"72",x"1e",x"66",x"c4"),
    46 => (x"87",x"f5",x"e9",x"49"),
    47 => (x"1e",x"4f",x"26",x"26"),
    48 => (x"bf",x"fe",x"cf",x"c2"),
    49 => (x"87",x"c8",x"e6",x"49"),
    50 => (x"48",x"ea",x"ef",x"c2"),
    51 => (x"c2",x"78",x"bf",x"e8"),
    52 => (x"ec",x"48",x"e6",x"ef"),
    53 => (x"ef",x"c2",x"78",x"bf"),
    54 => (x"49",x"4a",x"bf",x"ea"),
    55 => (x"ca",x"99",x"ff",x"cf"),
    56 => (x"48",x"72",x"2a",x"b7"),
    57 => (x"ef",x"c2",x"b0",x"71"),
    58 => (x"4f",x"26",x"58",x"f2"),
    59 => (x"5c",x"5b",x"5e",x"0e"),
    60 => (x"4b",x"71",x"0e",x"5d"),
    61 => (x"c2",x"87",x"c8",x"ff"),
    62 => (x"c0",x"48",x"e5",x"ef"),
    63 => (x"e5",x"49",x"73",x"50"),
    64 => (x"49",x"70",x"87",x"f5"),
    65 => (x"cb",x"9c",x"c2",x"4c"),
    66 => (x"f9",x"cb",x"49",x"ee"),
    67 => (x"4d",x"49",x"70",x"87"),
    68 => (x"97",x"e5",x"ef",x"c2"),
    69 => (x"e2",x"c1",x"05",x"bf"),
    70 => (x"49",x"66",x"d0",x"87"),
    71 => (x"bf",x"ee",x"ef",x"c2"),
    72 => (x"87",x"d6",x"05",x"99"),
    73 => (x"c2",x"49",x"66",x"d4"),
    74 => (x"99",x"bf",x"e6",x"ef"),
    75 => (x"73",x"87",x"cb",x"05"),
    76 => (x"87",x"c3",x"e5",x"49"),
    77 => (x"c1",x"02",x"98",x"70"),
    78 => (x"4c",x"c1",x"87",x"c1"),
    79 => (x"75",x"87",x"c0",x"fe"),
    80 => (x"87",x"ce",x"cb",x"49"),
    81 => (x"c6",x"02",x"98",x"70"),
    82 => (x"e5",x"ef",x"c2",x"87"),
    83 => (x"c2",x"50",x"c1",x"48"),
    84 => (x"bf",x"97",x"e5",x"ef"),
    85 => (x"87",x"e3",x"c0",x"05"),
    86 => (x"bf",x"ee",x"ef",x"c2"),
    87 => (x"99",x"66",x"d0",x"49"),
    88 => (x"87",x"d6",x"ff",x"05"),
    89 => (x"bf",x"e6",x"ef",x"c2"),
    90 => (x"99",x"66",x"d4",x"49"),
    91 => (x"87",x"ca",x"ff",x"05"),
    92 => (x"c2",x"e4",x"49",x"73"),
    93 => (x"05",x"98",x"70",x"87"),
    94 => (x"74",x"87",x"ff",x"fe"),
    95 => (x"87",x"dc",x"fb",x"48"),
    96 => (x"5c",x"5b",x"5e",x"0e"),
    97 => (x"86",x"f4",x"0e",x"5d"),
    98 => (x"ec",x"4c",x"4d",x"c0"),
    99 => (x"a6",x"c4",x"7e",x"bf"),
   100 => (x"f2",x"ef",x"c2",x"48"),
   101 => (x"1e",x"c1",x"78",x"bf"),
   102 => (x"49",x"c7",x"1e",x"c0"),
   103 => (x"c8",x"87",x"cd",x"fd"),
   104 => (x"02",x"98",x"70",x"86"),
   105 => (x"49",x"ff",x"87",x"cd"),
   106 => (x"c1",x"87",x"cc",x"fb"),
   107 => (x"c6",x"e3",x"49",x"da"),
   108 => (x"c2",x"4d",x"c1",x"87"),
   109 => (x"bf",x"97",x"e5",x"ef"),
   110 => (x"d5",x"87",x"c3",x"02"),
   111 => (x"ef",x"c2",x"87",x"de"),
   112 => (x"c2",x"4b",x"bf",x"ea"),
   113 => (x"05",x"bf",x"fe",x"cf"),
   114 => (x"c4",x"87",x"da",x"c1"),
   115 => (x"c0",x"c2",x"48",x"a6"),
   116 => (x"c2",x"78",x"c0",x"c0"),
   117 => (x"6e",x"7e",x"ee",x"dd"),
   118 => (x"6e",x"49",x"bf",x"97"),
   119 => (x"70",x"80",x"c1",x"48"),
   120 => (x"d2",x"e2",x"71",x"7e"),
   121 => (x"02",x"98",x"70",x"87"),
   122 => (x"66",x"c4",x"87",x"c3"),
   123 => (x"48",x"66",x"c4",x"b3"),
   124 => (x"c8",x"28",x"b7",x"c1"),
   125 => (x"98",x"70",x"58",x"a6"),
   126 => (x"87",x"db",x"ff",x"05"),
   127 => (x"e1",x"49",x"fd",x"c3"),
   128 => (x"fa",x"c3",x"87",x"f5"),
   129 => (x"87",x"ef",x"e1",x"49"),
   130 => (x"ff",x"cf",x"49",x"73"),
   131 => (x"c0",x"1e",x"71",x"99"),
   132 => (x"87",x"dd",x"fa",x"49"),
   133 => (x"b7",x"ca",x"49",x"73"),
   134 => (x"c1",x"1e",x"71",x"29"),
   135 => (x"87",x"d1",x"fa",x"49"),
   136 => (x"ff",x"c5",x"86",x"c8"),
   137 => (x"ee",x"ef",x"c2",x"87"),
   138 => (x"02",x"9b",x"4b",x"bf"),
   139 => (x"cf",x"c2",x"87",x"dd"),
   140 => (x"c7",x"49",x"bf",x"fa"),
   141 => (x"98",x"70",x"87",x"dc"),
   142 => (x"c0",x"87",x"c4",x"05"),
   143 => (x"c2",x"87",x"d2",x"4b"),
   144 => (x"c1",x"c7",x"49",x"e0"),
   145 => (x"fe",x"cf",x"c2",x"87"),
   146 => (x"c2",x"87",x"c6",x"58"),
   147 => (x"c0",x"48",x"fa",x"cf"),
   148 => (x"c2",x"49",x"73",x"78"),
   149 => (x"87",x"cd",x"05",x"99"),
   150 => (x"e0",x"49",x"eb",x"c3"),
   151 => (x"49",x"70",x"87",x"d9"),
   152 => (x"c2",x"02",x"99",x"c2"),
   153 => (x"73",x"4c",x"fb",x"87"),
   154 => (x"05",x"99",x"c1",x"49"),
   155 => (x"f4",x"c3",x"87",x"cd"),
   156 => (x"87",x"c3",x"e0",x"49"),
   157 => (x"99",x"c2",x"49",x"70"),
   158 => (x"fa",x"87",x"c2",x"02"),
   159 => (x"c8",x"49",x"73",x"4c"),
   160 => (x"87",x"ce",x"05",x"99"),
   161 => (x"ff",x"49",x"f5",x"c3"),
   162 => (x"70",x"87",x"ec",x"df"),
   163 => (x"02",x"99",x"c2",x"49"),
   164 => (x"ef",x"c2",x"87",x"d5"),
   165 => (x"ca",x"02",x"bf",x"f6"),
   166 => (x"88",x"c1",x"48",x"87"),
   167 => (x"58",x"fa",x"ef",x"c2"),
   168 => (x"ff",x"87",x"c2",x"c0"),
   169 => (x"73",x"4d",x"c1",x"4c"),
   170 => (x"05",x"99",x"c4",x"49"),
   171 => (x"f2",x"c3",x"87",x"ce"),
   172 => (x"c2",x"df",x"ff",x"49"),
   173 => (x"c2",x"49",x"70",x"87"),
   174 => (x"87",x"dc",x"02",x"99"),
   175 => (x"bf",x"f6",x"ef",x"c2"),
   176 => (x"b7",x"c7",x"48",x"7e"),
   177 => (x"cb",x"c0",x"03",x"a8"),
   178 => (x"c1",x"48",x"6e",x"87"),
   179 => (x"fa",x"ef",x"c2",x"80"),
   180 => (x"87",x"c2",x"c0",x"58"),
   181 => (x"4d",x"c1",x"4c",x"fe"),
   182 => (x"ff",x"49",x"fd",x"c3"),
   183 => (x"70",x"87",x"d8",x"de"),
   184 => (x"02",x"99",x"c2",x"49"),
   185 => (x"c2",x"87",x"d5",x"c0"),
   186 => (x"02",x"bf",x"f6",x"ef"),
   187 => (x"c2",x"87",x"c9",x"c0"),
   188 => (x"c0",x"48",x"f6",x"ef"),
   189 => (x"87",x"c2",x"c0",x"78"),
   190 => (x"4d",x"c1",x"4c",x"fd"),
   191 => (x"ff",x"49",x"fa",x"c3"),
   192 => (x"70",x"87",x"f4",x"dd"),
   193 => (x"02",x"99",x"c2",x"49"),
   194 => (x"c2",x"87",x"d9",x"c0"),
   195 => (x"48",x"bf",x"f6",x"ef"),
   196 => (x"03",x"a8",x"b7",x"c7"),
   197 => (x"c2",x"87",x"c9",x"c0"),
   198 => (x"c7",x"48",x"f6",x"ef"),
   199 => (x"87",x"c2",x"c0",x"78"),
   200 => (x"4d",x"c1",x"4c",x"fc"),
   201 => (x"03",x"ac",x"b7",x"c0"),
   202 => (x"c4",x"87",x"d1",x"c0"),
   203 => (x"d8",x"c1",x"4a",x"66"),
   204 => (x"c0",x"02",x"6a",x"82"),
   205 => (x"4b",x"6a",x"87",x"c6"),
   206 => (x"0f",x"73",x"49",x"74"),
   207 => (x"f0",x"c3",x"1e",x"c0"),
   208 => (x"49",x"da",x"c1",x"1e"),
   209 => (x"c8",x"87",x"e5",x"f6"),
   210 => (x"02",x"98",x"70",x"86"),
   211 => (x"c8",x"87",x"e2",x"c0"),
   212 => (x"ef",x"c2",x"48",x"a6"),
   213 => (x"c8",x"78",x"bf",x"f6"),
   214 => (x"91",x"cb",x"49",x"66"),
   215 => (x"71",x"48",x"66",x"c4"),
   216 => (x"6e",x"7e",x"70",x"80"),
   217 => (x"c8",x"c0",x"02",x"bf"),
   218 => (x"4b",x"bf",x"6e",x"87"),
   219 => (x"73",x"49",x"66",x"c8"),
   220 => (x"02",x"9d",x"75",x"0f"),
   221 => (x"c2",x"87",x"c8",x"c0"),
   222 => (x"49",x"bf",x"f6",x"ef"),
   223 => (x"c2",x"87",x"d3",x"f2"),
   224 => (x"02",x"bf",x"c2",x"d0"),
   225 => (x"49",x"87",x"dd",x"c0"),
   226 => (x"70",x"87",x"c7",x"c2"),
   227 => (x"d3",x"c0",x"02",x"98"),
   228 => (x"f6",x"ef",x"c2",x"87"),
   229 => (x"f9",x"f1",x"49",x"bf"),
   230 => (x"f3",x"49",x"c0",x"87"),
   231 => (x"d0",x"c2",x"87",x"d9"),
   232 => (x"78",x"c0",x"48",x"c2"),
   233 => (x"f3",x"f2",x"8e",x"f4"),
   234 => (x"5b",x"5e",x"0e",x"87"),
   235 => (x"1e",x"0e",x"5d",x"5c"),
   236 => (x"ef",x"c2",x"4c",x"71"),
   237 => (x"c1",x"49",x"bf",x"f2"),
   238 => (x"c1",x"4d",x"a1",x"cd"),
   239 => (x"7e",x"69",x"81",x"d1"),
   240 => (x"cf",x"02",x"9c",x"74"),
   241 => (x"4b",x"a5",x"c4",x"87"),
   242 => (x"ef",x"c2",x"7b",x"74"),
   243 => (x"f2",x"49",x"bf",x"f2"),
   244 => (x"7b",x"6e",x"87",x"d2"),
   245 => (x"c4",x"05",x"9c",x"74"),
   246 => (x"c2",x"4b",x"c0",x"87"),
   247 => (x"73",x"4b",x"c1",x"87"),
   248 => (x"87",x"d3",x"f2",x"49"),
   249 => (x"c7",x"02",x"66",x"d4"),
   250 => (x"87",x"da",x"49",x"87"),
   251 => (x"87",x"c2",x"4a",x"70"),
   252 => (x"d0",x"c2",x"4a",x"c0"),
   253 => (x"f1",x"26",x"5a",x"c6"),
   254 => (x"00",x"00",x"87",x"e2"),
   255 => (x"00",x"00",x"00",x"00"),
   256 => (x"00",x"00",x"00",x"00"),
   257 => (x"71",x"1e",x"00",x"00"),
   258 => (x"bf",x"c8",x"ff",x"4a"),
   259 => (x"48",x"a1",x"72",x"49"),
   260 => (x"ff",x"1e",x"4f",x"26"),
   261 => (x"fe",x"89",x"bf",x"c8"),
   262 => (x"c0",x"c0",x"c0",x"c0"),
   263 => (x"c4",x"01",x"a9",x"c0"),
   264 => (x"c2",x"4a",x"c0",x"87"),
   265 => (x"72",x"4a",x"c1",x"87"),
   266 => (x"0e",x"4f",x"26",x"48"),
   267 => (x"5d",x"5c",x"5b",x"5e"),
   268 => (x"ff",x"4b",x"71",x"0e"),
   269 => (x"66",x"d0",x"4c",x"d4"),
   270 => (x"d6",x"78",x"c0",x"48"),
   271 => (x"f6",x"da",x"ff",x"49"),
   272 => (x"7c",x"ff",x"c3",x"87"),
   273 => (x"ff",x"c3",x"49",x"6c"),
   274 => (x"49",x"4d",x"71",x"99"),
   275 => (x"c1",x"99",x"f0",x"c3"),
   276 => (x"cb",x"05",x"a9",x"e0"),
   277 => (x"7c",x"ff",x"c3",x"87"),
   278 => (x"98",x"c3",x"48",x"6c"),
   279 => (x"78",x"08",x"66",x"d0"),
   280 => (x"6c",x"7c",x"ff",x"c3"),
   281 => (x"31",x"c8",x"49",x"4a"),
   282 => (x"6c",x"7c",x"ff",x"c3"),
   283 => (x"72",x"b2",x"71",x"4a"),
   284 => (x"c3",x"31",x"c8",x"49"),
   285 => (x"4a",x"6c",x"7c",x"ff"),
   286 => (x"49",x"72",x"b2",x"71"),
   287 => (x"ff",x"c3",x"31",x"c8"),
   288 => (x"71",x"4a",x"6c",x"7c"),
   289 => (x"48",x"d0",x"ff",x"b2"),
   290 => (x"73",x"78",x"e0",x"c0"),
   291 => (x"87",x"c2",x"02",x"9b"),
   292 => (x"48",x"75",x"7b",x"72"),
   293 => (x"4c",x"26",x"4d",x"26"),
   294 => (x"4f",x"26",x"4b",x"26"),
   295 => (x"0e",x"4f",x"26",x"1e"),
   296 => (x"0e",x"5c",x"5b",x"5e"),
   297 => (x"1e",x"76",x"86",x"f8"),
   298 => (x"fd",x"49",x"a6",x"c8"),
   299 => (x"86",x"c4",x"87",x"fd"),
   300 => (x"48",x"6e",x"4b",x"70"),
   301 => (x"c2",x"01",x"a8",x"c0"),
   302 => (x"4a",x"73",x"87",x"f0"),
   303 => (x"c1",x"9a",x"f0",x"c3"),
   304 => (x"c7",x"02",x"aa",x"d0"),
   305 => (x"aa",x"e0",x"c1",x"87"),
   306 => (x"87",x"de",x"c2",x"05"),
   307 => (x"99",x"c8",x"49",x"73"),
   308 => (x"ff",x"87",x"c3",x"02"),
   309 => (x"4c",x"73",x"87",x"c6"),
   310 => (x"ac",x"c2",x"9c",x"c3"),
   311 => (x"87",x"c2",x"c1",x"05"),
   312 => (x"c9",x"49",x"66",x"c4"),
   313 => (x"c4",x"1e",x"71",x"31"),
   314 => (x"92",x"d4",x"4a",x"66"),
   315 => (x"49",x"fa",x"ef",x"c2"),
   316 => (x"d2",x"fe",x"81",x"72"),
   317 => (x"49",x"d8",x"87",x"f9"),
   318 => (x"87",x"fb",x"d7",x"ff"),
   319 => (x"c2",x"1e",x"c0",x"c8"),
   320 => (x"fd",x"49",x"ea",x"de"),
   321 => (x"ff",x"87",x"d4",x"ef"),
   322 => (x"e0",x"c0",x"48",x"d0"),
   323 => (x"ea",x"de",x"c2",x"78"),
   324 => (x"4a",x"66",x"cc",x"1e"),
   325 => (x"ef",x"c2",x"92",x"d4"),
   326 => (x"81",x"72",x"49",x"fa"),
   327 => (x"87",x"cc",x"d1",x"fe"),
   328 => (x"ac",x"c1",x"86",x"cc"),
   329 => (x"87",x"c2",x"c1",x"05"),
   330 => (x"c9",x"49",x"66",x"c4"),
   331 => (x"c4",x"1e",x"71",x"31"),
   332 => (x"92",x"d4",x"4a",x"66"),
   333 => (x"49",x"fa",x"ef",x"c2"),
   334 => (x"d1",x"fe",x"81",x"72"),
   335 => (x"de",x"c2",x"87",x"f1"),
   336 => (x"66",x"c8",x"1e",x"ea"),
   337 => (x"c2",x"92",x"d4",x"4a"),
   338 => (x"72",x"49",x"fa",x"ef"),
   339 => (x"d8",x"cf",x"fe",x"81"),
   340 => (x"ff",x"49",x"d7",x"87"),
   341 => (x"c8",x"87",x"e0",x"d6"),
   342 => (x"de",x"c2",x"1e",x"c0"),
   343 => (x"ed",x"fd",x"49",x"ea"),
   344 => (x"86",x"cc",x"87",x"e3"),
   345 => (x"c0",x"48",x"d0",x"ff"),
   346 => (x"8e",x"f8",x"78",x"e0"),
   347 => (x"0e",x"87",x"e7",x"fc"),
   348 => (x"5d",x"5c",x"5b",x"5e"),
   349 => (x"4d",x"71",x"1e",x"0e"),
   350 => (x"d4",x"4c",x"d4",x"ff"),
   351 => (x"c3",x"48",x"7e",x"66"),
   352 => (x"c5",x"06",x"a8",x"b7"),
   353 => (x"c1",x"48",x"c0",x"87"),
   354 => (x"49",x"75",x"87",x"e2"),
   355 => (x"87",x"f0",x"df",x"fe"),
   356 => (x"66",x"c4",x"1e",x"75"),
   357 => (x"c2",x"93",x"d4",x"4b"),
   358 => (x"73",x"83",x"fa",x"ef"),
   359 => (x"ec",x"ca",x"fe",x"49"),
   360 => (x"6b",x"83",x"c8",x"87"),
   361 => (x"48",x"d0",x"ff",x"4b"),
   362 => (x"dd",x"78",x"e1",x"c8"),
   363 => (x"c3",x"49",x"73",x"7c"),
   364 => (x"7c",x"71",x"99",x"ff"),
   365 => (x"b7",x"c8",x"49",x"73"),
   366 => (x"99",x"ff",x"c3",x"29"),
   367 => (x"49",x"73",x"7c",x"71"),
   368 => (x"c3",x"29",x"b7",x"d0"),
   369 => (x"7c",x"71",x"99",x"ff"),
   370 => (x"b7",x"d8",x"49",x"73"),
   371 => (x"c0",x"7c",x"71",x"29"),
   372 => (x"7c",x"7c",x"7c",x"7c"),
   373 => (x"7c",x"7c",x"7c",x"7c"),
   374 => (x"7c",x"7c",x"7c",x"7c"),
   375 => (x"c4",x"78",x"e0",x"c0"),
   376 => (x"49",x"dc",x"1e",x"66"),
   377 => (x"87",x"f4",x"d4",x"ff"),
   378 => (x"48",x"73",x"86",x"c8"),
   379 => (x"87",x"e4",x"fa",x"26"),
   380 => (x"5c",x"5b",x"5e",x"0e"),
   381 => (x"71",x"1e",x"0e",x"5d"),
   382 => (x"4b",x"d4",x"ff",x"7e"),
   383 => (x"f0",x"c2",x"1e",x"6e"),
   384 => (x"c9",x"fe",x"49",x"ce"),
   385 => (x"86",x"c4",x"87",x"c7"),
   386 => (x"02",x"9d",x"4d",x"70"),
   387 => (x"c2",x"87",x"c3",x"c3"),
   388 => (x"4c",x"bf",x"d6",x"f0"),
   389 => (x"dd",x"fe",x"49",x"6e"),
   390 => (x"d0",x"ff",x"87",x"e6"),
   391 => (x"78",x"c5",x"c8",x"48"),
   392 => (x"c0",x"7b",x"d6",x"c1"),
   393 => (x"c1",x"7b",x"15",x"4a"),
   394 => (x"b7",x"e0",x"c0",x"82"),
   395 => (x"87",x"f5",x"04",x"aa"),
   396 => (x"c4",x"48",x"d0",x"ff"),
   397 => (x"78",x"c5",x"c8",x"78"),
   398 => (x"c1",x"7b",x"d3",x"c1"),
   399 => (x"74",x"78",x"c4",x"7b"),
   400 => (x"fc",x"c1",x"02",x"9c"),
   401 => (x"ea",x"de",x"c2",x"87"),
   402 => (x"4d",x"c0",x"c8",x"7e"),
   403 => (x"ac",x"b7",x"c0",x"8c"),
   404 => (x"c8",x"87",x"c6",x"03"),
   405 => (x"c0",x"4d",x"a4",x"c0"),
   406 => (x"db",x"eb",x"c2",x"4c"),
   407 => (x"d0",x"49",x"bf",x"97"),
   408 => (x"87",x"d2",x"02",x"99"),
   409 => (x"f0",x"c2",x"1e",x"c0"),
   410 => (x"ca",x"fe",x"49",x"ce"),
   411 => (x"86",x"c4",x"87",x"fb"),
   412 => (x"c0",x"4a",x"49",x"70"),
   413 => (x"de",x"c2",x"87",x"ef"),
   414 => (x"f0",x"c2",x"1e",x"ea"),
   415 => (x"ca",x"fe",x"49",x"ce"),
   416 => (x"86",x"c4",x"87",x"e7"),
   417 => (x"ff",x"4a",x"49",x"70"),
   418 => (x"c5",x"c8",x"48",x"d0"),
   419 => (x"7b",x"d4",x"c1",x"78"),
   420 => (x"7b",x"bf",x"97",x"6e"),
   421 => (x"80",x"c1",x"48",x"6e"),
   422 => (x"8d",x"c1",x"7e",x"70"),
   423 => (x"87",x"f0",x"ff",x"05"),
   424 => (x"c4",x"48",x"d0",x"ff"),
   425 => (x"05",x"9a",x"72",x"78"),
   426 => (x"48",x"c0",x"87",x"c5"),
   427 => (x"c1",x"87",x"e5",x"c0"),
   428 => (x"ce",x"f0",x"c2",x"1e"),
   429 => (x"cf",x"c8",x"fe",x"49"),
   430 => (x"74",x"86",x"c4",x"87"),
   431 => (x"c4",x"fe",x"05",x"9c"),
   432 => (x"48",x"d0",x"ff",x"87"),
   433 => (x"c1",x"78",x"c5",x"c8"),
   434 => (x"7b",x"c0",x"7b",x"d3"),
   435 => (x"48",x"c1",x"78",x"c4"),
   436 => (x"48",x"c0",x"87",x"c2"),
   437 => (x"26",x"4d",x"26",x"26"),
   438 => (x"26",x"4b",x"26",x"4c"),
   439 => (x"5b",x"5e",x"0e",x"4f"),
   440 => (x"4b",x"71",x"0e",x"5c"),
   441 => (x"d8",x"02",x"66",x"cc"),
   442 => (x"f0",x"c0",x"4c",x"87"),
   443 => (x"87",x"d8",x"02",x"8c"),
   444 => (x"8a",x"c1",x"4a",x"74"),
   445 => (x"8a",x"87",x"d1",x"02"),
   446 => (x"8a",x"87",x"cd",x"02"),
   447 => (x"d7",x"87",x"c9",x"02"),
   448 => (x"fb",x"49",x"73",x"87"),
   449 => (x"87",x"d0",x"87",x"ea"),
   450 => (x"49",x"c0",x"1e",x"74"),
   451 => (x"74",x"87",x"e0",x"f9"),
   452 => (x"f9",x"49",x"73",x"1e"),
   453 => (x"86",x"c8",x"87",x"d9"),
   454 => (x"00",x"87",x"fc",x"fe"),
   455 => (x"ea",x"dd",x"c2",x"1e"),
   456 => (x"b9",x"c1",x"49",x"bf"),
   457 => (x"59",x"ee",x"dd",x"c2"),
   458 => (x"c3",x"48",x"d4",x"ff"),
   459 => (x"d0",x"ff",x"78",x"ff"),
   460 => (x"78",x"e1",x"c8",x"48"),
   461 => (x"c1",x"48",x"d4",x"ff"),
   462 => (x"71",x"31",x"c4",x"78"),
   463 => (x"48",x"d0",x"ff",x"78"),
   464 => (x"26",x"78",x"e0",x"c0"),
   465 => (x"dd",x"c2",x"1e",x"4f"),
   466 => (x"f0",x"c2",x"1e",x"de"),
   467 => (x"c3",x"fe",x"49",x"ce"),
   468 => (x"86",x"c4",x"87",x"fb"),
   469 => (x"c3",x"02",x"98",x"70"),
   470 => (x"87",x"c0",x"ff",x"87"),
   471 => (x"35",x"31",x"4f",x"26"),
   472 => (x"20",x"5a",x"48",x"4b"),
   473 => (x"46",x"43",x"20",x"20"),
   474 => (x"00",x"00",x"00",x"47"),
   475 => (x"9f",x"1a",x"00",x"00"),
   476 => (x"14",x"11",x"12",x"58"),
   477 => (x"23",x"1c",x"1b",x"1d"),
   478 => (x"59",x"5a",x"a7",x"4a"),
   479 => (x"f2",x"f5",x"94",x"91"),
   480 => (x"f2",x"f5",x"f4",x"eb"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

