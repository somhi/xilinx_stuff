library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom1 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"e4f0c287",
    12 => x"86c0c64e",
    13 => x"49e4f0c2",
    14 => x"48c4dec2",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087f8db",
    19 => x"1e87fc98",
    20 => x"1e731e72",
    21 => x"02114812",
    22 => x"c34b87ca",
    23 => x"739b98df",
    24 => x"87f00288",
    25 => x"4a264b26",
    26 => x"731e4f26",
    27 => x"c11e721e",
    28 => x"87ca048b",
    29 => x"02114812",
    30 => x"028887c4",
    31 => x"4a2687f1",
    32 => x"4f264b26",
    33 => x"731e741e",
    34 => x"c11e721e",
    35 => x"87d0048b",
    36 => x"02114812",
    37 => x"c34c87ca",
    38 => x"749c98df",
    39 => x"87eb0288",
    40 => x"4b264a26",
    41 => x"4f264c26",
    42 => x"8148731e",
    43 => x"c502a973",
    44 => x"05531287",
    45 => x"4f2687f6",
    46 => x"4a66c41e",
    47 => x"51124871",
    48 => x"2687fb05",
    49 => x"48111e4f",
    50 => x"7808d4ff",
    51 => x"c14866c4",
    52 => x"58a6c888",
    53 => x"ed059870",
    54 => x"1e4f2687",
    55 => x"c348d4ff",
    56 => x"516878ff",
    57 => x"c14866c4",
    58 => x"58a6c888",
    59 => x"eb059870",
    60 => x"1e4f2687",
    61 => x"d4ff1e73",
    62 => x"7bffc34b",
    63 => x"ffc34a6b",
    64 => x"c8496b7b",
    65 => x"c3b17232",
    66 => x"4a6b7bff",
    67 => x"b27131c8",
    68 => x"6b7bffc3",
    69 => x"7232c849",
    70 => x"c44871b1",
    71 => x"264d2687",
    72 => x"264b264c",
    73 => x"5b5e0e4f",
    74 => x"710e5d5c",
    75 => x"4cd4ff4a",
    76 => x"ffc34972",
    77 => x"c27c7199",
    78 => x"05bfc4de",
    79 => x"66d087c8",
    80 => x"d430c948",
    81 => x"66d058a6",
    82 => x"c329d849",
    83 => x"7c7199ff",
    84 => x"d04966d0",
    85 => x"99ffc329",
    86 => x"66d07c71",
    87 => x"c329c849",
    88 => x"7c7199ff",
    89 => x"c34966d0",
    90 => x"7c7199ff",
    91 => x"29d04972",
    92 => x"7199ffc3",
    93 => x"c94b6c7c",
    94 => x"c34dfff0",
    95 => x"d005abff",
    96 => x"7cffc387",
    97 => x"8dc14b6c",
    98 => x"c387c602",
    99 => x"f002abff",
   100 => x"fe487387",
   101 => x"c01e87c7",
   102 => x"48d4ff49",
   103 => x"c178ffc3",
   104 => x"b7c8c381",
   105 => x"87f104a9",
   106 => x"731e4f26",
   107 => x"c487e71e",
   108 => x"c04bdff8",
   109 => x"f0ffc01e",
   110 => x"fd49f7c1",
   111 => x"86c487e7",
   112 => x"c005a8c1",
   113 => x"d4ff87ea",
   114 => x"78ffc348",
   115 => x"c0c0c0c1",
   116 => x"c01ec0c0",
   117 => x"e9c1f0e1",
   118 => x"87c9fd49",
   119 => x"987086c4",
   120 => x"ff87ca05",
   121 => x"ffc348d4",
   122 => x"cb48c178",
   123 => x"87e6fe87",
   124 => x"fe058bc1",
   125 => x"48c087fd",
   126 => x"1e87e6fc",
   127 => x"d4ff1e73",
   128 => x"78ffc348",
   129 => x"1ec04bd3",
   130 => x"c1f0ffc0",
   131 => x"d4fc49c1",
   132 => x"7086c487",
   133 => x"87ca0598",
   134 => x"c348d4ff",
   135 => x"48c178ff",
   136 => x"f1fd87cb",
   137 => x"058bc187",
   138 => x"c087dbff",
   139 => x"87f1fb48",
   140 => x"5c5b5e0e",
   141 => x"4cd4ff0e",
   142 => x"c687dbfd",
   143 => x"e1c01eea",
   144 => x"49c8c1f0",
   145 => x"c487defb",
   146 => x"02a8c186",
   147 => x"eafe87c8",
   148 => x"c148c087",
   149 => x"dafa87e2",
   150 => x"cf497087",
   151 => x"c699ffff",
   152 => x"c802a9ea",
   153 => x"87d3fe87",
   154 => x"cbc148c0",
   155 => x"7cffc387",
   156 => x"fc4bf1c0",
   157 => x"987087f4",
   158 => x"87ebc002",
   159 => x"ffc01ec0",
   160 => x"49fac1f0",
   161 => x"c487defa",
   162 => x"05987086",
   163 => x"ffc387d9",
   164 => x"c3496c7c",
   165 => x"7c7c7cff",
   166 => x"99c0c17c",
   167 => x"c187c402",
   168 => x"c087d548",
   169 => x"c287d148",
   170 => x"87c405ab",
   171 => x"87c848c0",
   172 => x"fe058bc1",
   173 => x"48c087fd",
   174 => x"1e87e4f9",
   175 => x"dec21e73",
   176 => x"78c148c4",
   177 => x"d0ff4bc7",
   178 => x"fb78c248",
   179 => x"d0ff87c8",
   180 => x"c078c348",
   181 => x"d0e5c01e",
   182 => x"f949c0c1",
   183 => x"86c487c7",
   184 => x"c105a8c1",
   185 => x"abc24b87",
   186 => x"c087c505",
   187 => x"87f9c048",
   188 => x"ff058bc1",
   189 => x"f7fc87d0",
   190 => x"c8dec287",
   191 => x"05987058",
   192 => x"1ec187cd",
   193 => x"c1f0ffc0",
   194 => x"d8f849d0",
   195 => x"ff86c487",
   196 => x"ffc348d4",
   197 => x"87e0c478",
   198 => x"58ccdec2",
   199 => x"c248d0ff",
   200 => x"48d4ff78",
   201 => x"c178ffc3",
   202 => x"87f5f748",
   203 => x"5c5b5e0e",
   204 => x"4a710e5d",
   205 => x"ff4dffc3",
   206 => x"7c754cd4",
   207 => x"c448d0ff",
   208 => x"7c7578c3",
   209 => x"ffc01e72",
   210 => x"49d8c1f0",
   211 => x"c487d6f7",
   212 => x"02987086",
   213 => x"48c087c5",
   214 => x"7587f0c0",
   215 => x"7cfec37c",
   216 => x"d41ec0c8",
   217 => x"dcf54966",
   218 => x"7586c487",
   219 => x"757c757c",
   220 => x"e0dad87c",
   221 => x"6c7c754b",
   222 => x"c5059949",
   223 => x"058bc187",
   224 => x"7c7587f3",
   225 => x"c248d0ff",
   226 => x"f648c178",
   227 => x"ff1e87cf",
   228 => x"d0ff4ad4",
   229 => x"78d1c448",
   230 => x"c17affc3",
   231 => x"87f80589",
   232 => x"731e4f26",
   233 => x"c54b711e",
   234 => x"4adfcdee",
   235 => x"c348d4ff",
   236 => x"486878ff",
   237 => x"02a8fec3",
   238 => x"8ac187c5",
   239 => x"7287ed05",
   240 => x"87c5059a",
   241 => x"eac048c0",
   242 => x"029b7387",
   243 => x"66c887cc",
   244 => x"f449731e",
   245 => x"86c487c5",
   246 => x"66c887c6",
   247 => x"87eefe49",
   248 => x"c348d4ff",
   249 => x"737878ff",
   250 => x"87c5059b",
   251 => x"d048d0ff",
   252 => x"f448c178",
   253 => x"731e87eb",
   254 => x"c04a711e",
   255 => x"48d4ff4b",
   256 => x"ff78ffc3",
   257 => x"c3c448d0",
   258 => x"48d4ff78",
   259 => x"7278ffc3",
   260 => x"f0ffc01e",
   261 => x"f449d1c1",
   262 => x"86c487cb",
   263 => x"cd059870",
   264 => x"1ec0c887",
   265 => x"fd4966cc",
   266 => x"86c487f8",
   267 => x"d0ff4b70",
   268 => x"7378c248",
   269 => x"87e9f348",
   270 => x"5c5b5e0e",
   271 => x"1ec00e5d",
   272 => x"c1f0ffc0",
   273 => x"dcf349c9",
   274 => x"c21ed287",
   275 => x"fd49ccde",
   276 => x"86c887d0",
   277 => x"84c14cc0",
   278 => x"04acb7d2",
   279 => x"dec287f8",
   280 => x"49bf97cc",
   281 => x"c199c0c3",
   282 => x"c005a9c0",
   283 => x"dec287e7",
   284 => x"49bf97d3",
   285 => x"dec231d0",
   286 => x"4abf97d4",
   287 => x"b17232c8",
   288 => x"97d5dec2",
   289 => x"71b14abf",
   290 => x"ffffcf4c",
   291 => x"84c19cff",
   292 => x"e7c134ca",
   293 => x"d5dec287",
   294 => x"c149bf97",
   295 => x"c299c631",
   296 => x"bf97d6de",
   297 => x"2ab7c74a",
   298 => x"dec2b172",
   299 => x"4abf97d1",
   300 => x"c29dcf4d",
   301 => x"bf97d2de",
   302 => x"ca9ac34a",
   303 => x"d3dec232",
   304 => x"c24bbf97",
   305 => x"c2b27333",
   306 => x"bf97d4de",
   307 => x"9bc0c34b",
   308 => x"732bb7c6",
   309 => x"c181c2b2",
   310 => x"70307148",
   311 => x"7548c149",
   312 => x"724d7030",
   313 => x"7184c14c",
   314 => x"b7c0c894",
   315 => x"87cc06ad",
   316 => x"2db734c1",
   317 => x"adb7c0c8",
   318 => x"87f4ff01",
   319 => x"dcf04874",
   320 => x"5b5e0e87",
   321 => x"f80e5d5c",
   322 => x"f2e6c286",
   323 => x"c278c048",
   324 => x"c01eeade",
   325 => x"87defb49",
   326 => x"987086c4",
   327 => x"c087c505",
   328 => x"87cec948",
   329 => x"7ec14dc0",
   330 => x"bfcbf2c0",
   331 => x"e0dfc249",
   332 => x"4bc8714a",
   333 => x"7087f3ec",
   334 => x"87c20598",
   335 => x"f2c07ec0",
   336 => x"c249bfc7",
   337 => x"714afcdf",
   338 => x"ddec4bc8",
   339 => x"05987087",
   340 => x"7ec087c2",
   341 => x"fdc0026e",
   342 => x"f0e5c287",
   343 => x"e6c24dbf",
   344 => x"7ebf9fe8",
   345 => x"ead6c548",
   346 => x"87c705a8",
   347 => x"bff0e5c2",
   348 => x"6e87ce4d",
   349 => x"d5e9ca48",
   350 => x"87c502a8",
   351 => x"f1c748c0",
   352 => x"eadec287",
   353 => x"f949751e",
   354 => x"86c487ec",
   355 => x"c5059870",
   356 => x"c748c087",
   357 => x"f2c087dc",
   358 => x"c249bfc7",
   359 => x"714afcdf",
   360 => x"c5eb4bc8",
   361 => x"05987087",
   362 => x"e6c287c8",
   363 => x"78c148f2",
   364 => x"f2c087da",
   365 => x"c249bfcb",
   366 => x"714ae0df",
   367 => x"e9ea4bc8",
   368 => x"02987087",
   369 => x"c087c5c0",
   370 => x"87e6c648",
   371 => x"97e8e6c2",
   372 => x"d5c149bf",
   373 => x"cdc005a9",
   374 => x"e9e6c287",
   375 => x"c249bf97",
   376 => x"c002a9ea",
   377 => x"48c087c5",
   378 => x"c287c7c6",
   379 => x"bf97eade",
   380 => x"e9c3487e",
   381 => x"cec002a8",
   382 => x"c3486e87",
   383 => x"c002a8eb",
   384 => x"48c087c5",
   385 => x"c287ebc5",
   386 => x"bf97f5de",
   387 => x"c0059949",
   388 => x"dec287cc",
   389 => x"49bf97f6",
   390 => x"c002a9c2",
   391 => x"48c087c5",
   392 => x"c287cfc5",
   393 => x"bf97f7de",
   394 => x"eee6c248",
   395 => x"484c7058",
   396 => x"e6c288c1",
   397 => x"dec258f2",
   398 => x"49bf97f8",
   399 => x"dec28175",
   400 => x"4abf97f9",
   401 => x"a17232c8",
   402 => x"ffeac27e",
   403 => x"c2786e48",
   404 => x"bf97fade",
   405 => x"58a6c848",
   406 => x"bff2e6c2",
   407 => x"87d4c202",
   408 => x"bfc7f2c0",
   409 => x"fcdfc249",
   410 => x"4bc8714a",
   411 => x"7087fbe7",
   412 => x"c5c00298",
   413 => x"c348c087",
   414 => x"e6c287f8",
   415 => x"c24cbfea",
   416 => x"c25cd3eb",
   417 => x"bf97cfdf",
   418 => x"c231c849",
   419 => x"bf97cedf",
   420 => x"c249a14a",
   421 => x"bf97d0df",
   422 => x"7232d04a",
   423 => x"dfc249a1",
   424 => x"4abf97d1",
   425 => x"a17232d8",
   426 => x"9166c449",
   427 => x"bfffeac2",
   428 => x"c7ebc281",
   429 => x"d7dfc259",
   430 => x"c84abf97",
   431 => x"d6dfc232",
   432 => x"a24bbf97",
   433 => x"d8dfc24a",
   434 => x"d04bbf97",
   435 => x"4aa27333",
   436 => x"97d9dfc2",
   437 => x"9bcf4bbf",
   438 => x"a27333d8",
   439 => x"cbebc24a",
   440 => x"c7ebc25a",
   441 => x"8ac24abf",
   442 => x"ebc29274",
   443 => x"a17248cb",
   444 => x"87cac178",
   445 => x"97fcdec2",
   446 => x"31c849bf",
   447 => x"97fbdec2",
   448 => x"49a14abf",
   449 => x"59fae6c2",
   450 => x"bff6e6c2",
   451 => x"c731c549",
   452 => x"29c981ff",
   453 => x"59d3ebc2",
   454 => x"97c1dfc2",
   455 => x"32c84abf",
   456 => x"97c0dfc2",
   457 => x"4aa24bbf",
   458 => x"6e9266c4",
   459 => x"cfebc282",
   460 => x"c7ebc25a",
   461 => x"c278c048",
   462 => x"7248c3eb",
   463 => x"ebc278a1",
   464 => x"ebc248d3",
   465 => x"c278bfc7",
   466 => x"c248d7eb",
   467 => x"78bfcbeb",
   468 => x"bff2e6c2",
   469 => x"87c9c002",
   470 => x"30c44874",
   471 => x"c9c07e70",
   472 => x"cfebc287",
   473 => x"30c448bf",
   474 => x"e6c27e70",
   475 => x"786e48f6",
   476 => x"8ef848c1",
   477 => x"4c264d26",
   478 => x"4f264b26",
   479 => x"5c5b5e0e",
   480 => x"4a710e5d",
   481 => x"bff2e6c2",
   482 => x"7287cb02",
   483 => x"722bc74b",
   484 => x"9cffc14c",
   485 => x"4b7287c9",
   486 => x"4c722bc8",
   487 => x"c29cffc3",
   488 => x"83bfffea",
   489 => x"bfc3f2c0",
   490 => x"87d902ab",
   491 => x"5bc7f2c0",
   492 => x"1eeadec2",
   493 => x"fdf04973",
   494 => x"7086c487",
   495 => x"87c50598",
   496 => x"e6c048c0",
   497 => x"f2e6c287",
   498 => x"87d202bf",
   499 => x"91c44974",
   500 => x"81eadec2",
   501 => x"ffcf4d69",
   502 => x"9dffffff",
   503 => x"497487cb",
   504 => x"dec291c2",
   505 => x"699f81ea",
   506 => x"fe48754d",
   507 => x"5e0e87c6",
   508 => x"0e5d5c5b",
   509 => x"c04d711e",
   510 => x"ca49c11e",
   511 => x"86c487ee",
   512 => x"029c4c70",
   513 => x"c287c0c1",
   514 => x"754afae6",
   515 => x"87ffe049",
   516 => x"c0029870",
   517 => x"4a7487f1",
   518 => x"4bcb4975",
   519 => x"7087e5e1",
   520 => x"e2c00298",
   521 => x"741ec087",
   522 => x"87c7029c",
   523 => x"c048a6c4",
   524 => x"c487c578",
   525 => x"78c148a6",
   526 => x"c94966c4",
   527 => x"86c487ee",
   528 => x"059c4c70",
   529 => x"7487c0ff",
   530 => x"e7fc2648",
   531 => x"5b5e0e87",
   532 => x"1e0e5d5c",
   533 => x"059b4b71",
   534 => x"48c087c5",
   535 => x"c887e5c1",
   536 => x"7dc04da3",
   537 => x"c70266d4",
   538 => x"9766d487",
   539 => x"87c505bf",
   540 => x"cfc148c0",
   541 => x"4966d487",
   542 => x"7087f3fd",
   543 => x"c1029c4c",
   544 => x"a4dc87c0",
   545 => x"da7d6949",
   546 => x"a3c449a4",
   547 => x"7a699f4a",
   548 => x"bff2e6c2",
   549 => x"d487d202",
   550 => x"699f49a4",
   551 => x"ffffc049",
   552 => x"d0487199",
   553 => x"c27e7030",
   554 => x"6e7ec087",
   555 => x"806a4849",
   556 => x"7bc07a70",
   557 => x"6a49a3cc",
   558 => x"49a3d079",
   559 => x"487479c0",
   560 => x"48c087c2",
   561 => x"87ecfa26",
   562 => x"5c5b5e0e",
   563 => x"4c710e5d",
   564 => x"48c3f2c0",
   565 => x"9c7478ff",
   566 => x"87cac102",
   567 => x"6949a4c8",
   568 => x"87c2c102",
   569 => x"6c4a66d0",
   570 => x"a6d48249",
   571 => x"4d66d05a",
   572 => x"eee6c2b9",
   573 => x"baff4abf",
   574 => x"99719972",
   575 => x"87e4c002",
   576 => x"6b4ba4c4",
   577 => x"87f4f949",
   578 => x"e6c27b70",
   579 => x"6c49bfea",
   580 => x"757c7181",
   581 => x"eee6c2b9",
   582 => x"baff4abf",
   583 => x"99719972",
   584 => x"87dcff05",
   585 => x"cbf97c75",
   586 => x"1e731e87",
   587 => x"029b4b71",
   588 => x"a3c887c7",
   589 => x"c5056949",
   590 => x"c048c087",
   591 => x"ebc287eb",
   592 => x"c44abfc3",
   593 => x"496949a3",
   594 => x"e6c289c2",
   595 => x"7191bfea",
   596 => x"e6c24aa2",
   597 => x"6b49bfee",
   598 => x"4aa27199",
   599 => x"721e66c8",
   600 => x"87d2ea49",
   601 => x"497086c4",
   602 => x"87ccf848",
   603 => x"711e731e",
   604 => x"c7029b4b",
   605 => x"49a3c887",
   606 => x"87c50569",
   607 => x"ebc048c0",
   608 => x"c3ebc287",
   609 => x"a3c44abf",
   610 => x"c2496949",
   611 => x"eae6c289",
   612 => x"a27191bf",
   613 => x"eee6c24a",
   614 => x"996b49bf",
   615 => x"c84aa271",
   616 => x"49721e66",
   617 => x"c487c5e6",
   618 => x"48497086",
   619 => x"0e87c9f7",
   620 => x"5d5c5b5e",
   621 => x"4b711e0e",
   622 => x"c94c66d4",
   623 => x"029b732c",
   624 => x"c887cfc1",
   625 => x"026949a3",
   626 => x"d087c7c1",
   627 => x"66d44da3",
   628 => x"eee6c27d",
   629 => x"b9ff49bf",
   630 => x"7e994a6b",
   631 => x"cd03ac71",
   632 => x"7d7bc087",
   633 => x"c44aa3cc",
   634 => x"796a49a3",
   635 => x"8c7287c2",
   636 => x"dd029c74",
   637 => x"731e4987",
   638 => x"87ccfb49",
   639 => x"66d486c4",
   640 => x"99ffc749",
   641 => x"c287cb02",
   642 => x"731eeade",
   643 => x"87d9fc49",
   644 => x"f52686c4",
   645 => x"731e87de",
   646 => x"9b4b711e",
   647 => x"87e4c002",
   648 => x"5bd7ebc2",
   649 => x"8ac24a73",
   650 => x"bfeae6c2",
   651 => x"ebc29249",
   652 => x"7248bfc3",
   653 => x"dbebc280",
   654 => x"c4487158",
   655 => x"fae6c230",
   656 => x"87edc058",
   657 => x"48d3ebc2",
   658 => x"bfc7ebc2",
   659 => x"d7ebc278",
   660 => x"cbebc248",
   661 => x"e6c278bf",
   662 => x"c902bff2",
   663 => x"eae6c287",
   664 => x"31c449bf",
   665 => x"ebc287c7",
   666 => x"c449bfcf",
   667 => x"fae6c231",
   668 => x"87c4f459",
   669 => x"5c5b5e0e",
   670 => x"c04a710e",
   671 => x"029a724b",
   672 => x"da87e1c0",
   673 => x"699f49a2",
   674 => x"f2e6c24b",
   675 => x"87cf02bf",
   676 => x"9f49a2d4",
   677 => x"c04c4969",
   678 => x"d09cffff",
   679 => x"c087c234",
   680 => x"b349744c",
   681 => x"edfd4973",
   682 => x"87caf387",
   683 => x"5c5b5e0e",
   684 => x"86f40e5d",
   685 => x"7ec04a71",
   686 => x"d8029a72",
   687 => x"e6dec287",
   688 => x"c278c048",
   689 => x"c248dede",
   690 => x"78bfd7eb",
   691 => x"48e2dec2",
   692 => x"bfd3ebc2",
   693 => x"c7e7c278",
   694 => x"c250c048",
   695 => x"49bff6e6",
   696 => x"bfe6dec2",
   697 => x"03aa714a",
   698 => x"7287ffc3",
   699 => x"0599cf49",
   700 => x"c287e0c0",
   701 => x"c21eeade",
   702 => x"49bfdede",
   703 => x"48dedec2",
   704 => x"7178a1c1",
   705 => x"c487efe3",
   706 => x"fff1c086",
   707 => x"eadec248",
   708 => x"c087cc78",
   709 => x"48bffff1",
   710 => x"c080e0c0",
   711 => x"c258c3f2",
   712 => x"48bfe6de",
   713 => x"dec280c1",
   714 => x"7f2758ea",
   715 => x"bf00000c",
   716 => x"9d4dbf97",
   717 => x"87e2c202",
   718 => x"02ade5c3",
   719 => x"c087dbc2",
   720 => x"4bbffff1",
   721 => x"1149a3cb",
   722 => x"05accf4c",
   723 => x"7587d2c1",
   724 => x"c199df49",
   725 => x"c291cd89",
   726 => x"c181fae6",
   727 => x"51124aa3",
   728 => x"124aa3c3",
   729 => x"4aa3c551",
   730 => x"a3c75112",
   731 => x"c951124a",
   732 => x"51124aa3",
   733 => x"124aa3ce",
   734 => x"4aa3d051",
   735 => x"a3d25112",
   736 => x"d451124a",
   737 => x"51124aa3",
   738 => x"124aa3d6",
   739 => x"4aa3d851",
   740 => x"a3dc5112",
   741 => x"de51124a",
   742 => x"51124aa3",
   743 => x"f9c07ec1",
   744 => x"c8497487",
   745 => x"eac00599",
   746 => x"d0497487",
   747 => x"87d00599",
   748 => x"c00266dc",
   749 => x"497387ca",
   750 => x"700f66dc",
   751 => x"87d30298",
   752 => x"c6c0056e",
   753 => x"fae6c287",
   754 => x"c050c048",
   755 => x"48bffff1",
   756 => x"c287e7c2",
   757 => x"c048c7e7",
   758 => x"e6c27e50",
   759 => x"c249bff6",
   760 => x"4abfe6de",
   761 => x"fc04aa71",
   762 => x"ebc287c1",
   763 => x"c005bfd7",
   764 => x"e6c287c8",
   765 => x"c102bff2",
   766 => x"f2c087fe",
   767 => x"78ff48c3",
   768 => x"bfe2dec2",
   769 => x"87f4ed49",
   770 => x"dec24970",
   771 => x"a6c459e6",
   772 => x"e2dec248",
   773 => x"e6c278bf",
   774 => x"c002bff2",
   775 => x"66c487d8",
   776 => x"ffffcf49",
   777 => x"a999f8ff",
   778 => x"87c5c002",
   779 => x"e1c04dc0",
   780 => x"c04dc187",
   781 => x"66c487dc",
   782 => x"f8ffcf49",
   783 => x"c002a999",
   784 => x"a6c887c8",
   785 => x"c078c048",
   786 => x"a6c887c5",
   787 => x"c878c148",
   788 => x"9d754d66",
   789 => x"87e0c005",
   790 => x"c24966c4",
   791 => x"eae6c289",
   792 => x"c2914abf",
   793 => x"4abfc3eb",
   794 => x"48dedec2",
   795 => x"c278a172",
   796 => x"c048e6de",
   797 => x"87e3f978",
   798 => x"8ef448c0",
   799 => x"0087f5eb",
   800 => x"ff000000",
   801 => x"8fffffff",
   802 => x"9800000c",
   803 => x"4600000c",
   804 => x"32335441",
   805 => x"00202020",
   806 => x"31544146",
   807 => x"20202036",
   808 => x"d4ff1e00",
   809 => x"78ffc348",
   810 => x"4f264868",
   811 => x"48d4ff1e",
   812 => x"ff78ffc3",
   813 => x"e1c848d0",
   814 => x"48d4ff78",
   815 => x"ebc278d4",
   816 => x"d4ff48db",
   817 => x"4f2650bf",
   818 => x"48d0ff1e",
   819 => x"2678e0c0",
   820 => x"ccff1e4f",
   821 => x"99497087",
   822 => x"c087c602",
   823 => x"f105a9fb",
   824 => x"26487187",
   825 => x"5b5e0e4f",
   826 => x"4b710e5c",
   827 => x"f0fe4cc0",
   828 => x"99497087",
   829 => x"87f9c002",
   830 => x"02a9ecc0",
   831 => x"c087f2c0",
   832 => x"c002a9fb",
   833 => x"66cc87eb",
   834 => x"c703acb7",
   835 => x"0266d087",
   836 => x"537187c2",
   837 => x"c2029971",
   838 => x"fe84c187",
   839 => x"497087c3",
   840 => x"87cd0299",
   841 => x"02a9ecc0",
   842 => x"fbc087c7",
   843 => x"d5ff05a9",
   844 => x"0266d087",
   845 => x"97c087c3",
   846 => x"a9ecc07b",
   847 => x"7487c405",
   848 => x"7487c54a",
   849 => x"8a0ac04a",
   850 => x"87c24872",
   851 => x"4c264d26",
   852 => x"4f264b26",
   853 => x"87c9fd1e",
   854 => x"f0c04970",
   855 => x"ca04a9b7",
   856 => x"b7f9c087",
   857 => x"87c301a9",
   858 => x"c189f0c0",
   859 => x"04a9b7c1",
   860 => x"dac187ca",
   861 => x"c301a9b7",
   862 => x"89f7c087",
   863 => x"4f264871",
   864 => x"5c5b5e0e",
   865 => x"ff4a710e",
   866 => x"49724cd4",
   867 => x"7087eac0",
   868 => x"c2029b4b",
   869 => x"ff8bc187",
   870 => x"c5c848d0",
   871 => x"7cd5c178",
   872 => x"31c64973",
   873 => x"97dbdcc2",
   874 => x"71484abf",
   875 => x"ff7c70b0",
   876 => x"78c448d0",
   877 => x"d5fe4873",
   878 => x"5b5e0e87",
   879 => x"f80e5d5c",
   880 => x"c04c7186",
   881 => x"87e4fb7e",
   882 => x"f9c04bc0",
   883 => x"49bf97e6",
   884 => x"cf04a9c0",
   885 => x"87f9fb87",
   886 => x"f9c083c1",
   887 => x"49bf97e6",
   888 => x"87f106ab",
   889 => x"97e6f9c0",
   890 => x"87cf02bf",
   891 => x"7087f2fa",
   892 => x"c6029949",
   893 => x"a9ecc087",
   894 => x"c087f105",
   895 => x"87e1fa4b",
   896 => x"dcfa4d70",
   897 => x"58a6c887",
   898 => x"7087d6fa",
   899 => x"c883c14a",
   900 => x"699749a4",
   901 => x"c702ad49",
   902 => x"adffc087",
   903 => x"87e7c005",
   904 => x"9749a4c9",
   905 => x"66c44969",
   906 => x"87c702a9",
   907 => x"a8ffc048",
   908 => x"ca87d405",
   909 => x"699749a4",
   910 => x"c602aa49",
   911 => x"aaffc087",
   912 => x"c187c405",
   913 => x"c087d07e",
   914 => x"c602adec",
   915 => x"adfbc087",
   916 => x"c087c405",
   917 => x"6e7ec14b",
   918 => x"87e1fe02",
   919 => x"7387e9f9",
   920 => x"fb8ef848",
   921 => x"0e0087e6",
   922 => x"5d5c5b5e",
   923 => x"4b711e0e",
   924 => x"ab4d4cc0",
   925 => x"87e8c004",
   926 => x"1ef9f6c0",
   927 => x"c4029d75",
   928 => x"c24ac087",
   929 => x"724ac187",
   930 => x"87e0f049",
   931 => x"7e7086c4",
   932 => x"056e84c1",
   933 => x"4c7387c2",
   934 => x"ac7385c1",
   935 => x"87d8ff06",
   936 => x"2626486e",
   937 => x"264c264d",
   938 => x"0e4f264b",
   939 => x"5d5c5b5e",
   940 => x"4c711e0e",
   941 => x"c291de49",
   942 => x"714df5eb",
   943 => x"026d9785",
   944 => x"c287ddc1",
   945 => x"4abfe0eb",
   946 => x"49728274",
   947 => x"7087d8fe",
   948 => x"c0026e7e",
   949 => x"ebc287f3",
   950 => x"4a6e4be8",
   951 => x"c7ff49cb",
   952 => x"4b7487c6",
   953 => x"ddc193cb",
   954 => x"83c483e7",
   955 => x"7be4fcc0",
   956 => x"c4c14974",
   957 => x"7b7587dc",
   958 => x"97f4ebc2",
   959 => x"c21e49bf",
   960 => x"c149e8eb",
   961 => x"c487d6df",
   962 => x"c1497486",
   963 => x"c087c3c4",
   964 => x"e2c5c149",
   965 => x"dcebc287",
   966 => x"c178c048",
   967 => x"87f9dc49",
   968 => x"87fffd26",
   969 => x"64616f4c",
   970 => x"2e676e69",
   971 => x"0e002e2e",
   972 => x"0e5c5b5e",
   973 => x"c24a4b71",
   974 => x"82bfe0eb",
   975 => x"e6fc4972",
   976 => x"9c4c7087",
   977 => x"4987c402",
   978 => x"c287e9ec",
   979 => x"c048e0eb",
   980 => x"dc49c178",
   981 => x"ccfd87c3",
   982 => x"5b5e0e87",
   983 => x"f40e5d5c",
   984 => x"eadec286",
   985 => x"c44cc04d",
   986 => x"78c048a6",
   987 => x"bfe0ebc2",
   988 => x"06a9c049",
   989 => x"c287c1c1",
   990 => x"9848eade",
   991 => x"87f8c002",
   992 => x"1ef9f6c0",
   993 => x"c70266c8",
   994 => x"48a6c487",
   995 => x"87c578c0",
   996 => x"c148a6c4",
   997 => x"4966c478",
   998 => x"c487d1ec",
   999 => x"c14d7086",
  1000 => x"4866c484",
  1001 => x"a6c880c1",
  1002 => x"e0ebc258",
  1003 => x"03ac49bf",
  1004 => x"9d7587c6",
  1005 => x"87c8ff05",
  1006 => x"9d754cc0",
  1007 => x"87e0c302",
  1008 => x"1ef9f6c0",
  1009 => x"c70266c8",
  1010 => x"48a6cc87",
  1011 => x"87c578c0",
  1012 => x"c148a6cc",
  1013 => x"4966cc78",
  1014 => x"c487d1eb",
  1015 => x"6e7e7086",
  1016 => x"87e9c202",
  1017 => x"81cb496e",
  1018 => x"d0496997",
  1019 => x"d6c10299",
  1020 => x"effcc087",
  1021 => x"cb49744a",
  1022 => x"e7ddc191",
  1023 => x"c8797281",
  1024 => x"51ffc381",
  1025 => x"91de4974",
  1026 => x"4df5ebc2",
  1027 => x"c1c28571",
  1028 => x"a5c17d97",
  1029 => x"51e0c049",
  1030 => x"97fae6c2",
  1031 => x"87d202bf",
  1032 => x"a5c284c1",
  1033 => x"fae6c24b",
  1034 => x"ff49db4a",
  1035 => x"c187f9c1",
  1036 => x"a5cd87db",
  1037 => x"c151c049",
  1038 => x"4ba5c284",
  1039 => x"49cb4a6e",
  1040 => x"87e4c1ff",
  1041 => x"c087c6c1",
  1042 => x"744aebfa",
  1043 => x"c191cb49",
  1044 => x"7281e7dd",
  1045 => x"fae6c279",
  1046 => x"d802bf97",
  1047 => x"de497487",
  1048 => x"c284c191",
  1049 => x"714bf5eb",
  1050 => x"fae6c283",
  1051 => x"ff49dd4a",
  1052 => x"d887f5c0",
  1053 => x"de4b7487",
  1054 => x"f5ebc293",
  1055 => x"49a3cb83",
  1056 => x"84c151c0",
  1057 => x"cb4a6e73",
  1058 => x"dbc0ff49",
  1059 => x"4866c487",
  1060 => x"a6c880c1",
  1061 => x"03acc758",
  1062 => x"6e87c5c0",
  1063 => x"87e0fc05",
  1064 => x"8ef44874",
  1065 => x"1e87fcf7",
  1066 => x"4b711e73",
  1067 => x"c191cb49",
  1068 => x"c881e7dd",
  1069 => x"dcc24aa1",
  1070 => x"501248db",
  1071 => x"c04aa1c9",
  1072 => x"1248e6f9",
  1073 => x"c281ca50",
  1074 => x"1148f4eb",
  1075 => x"f4ebc250",
  1076 => x"1e49bf97",
  1077 => x"d8c149c0",
  1078 => x"ebc287c3",
  1079 => x"78de48dc",
  1080 => x"f4d549c1",
  1081 => x"fef62687",
  1082 => x"4a711e87",
  1083 => x"c191cb49",
  1084 => x"c881e7dd",
  1085 => x"c2481181",
  1086 => x"c258e0eb",
  1087 => x"c048e0eb",
  1088 => x"d549c178",
  1089 => x"4f2687d3",
  1090 => x"c049c01e",
  1091 => x"2687e8fd",
  1092 => x"99711e4f",
  1093 => x"c187d202",
  1094 => x"c048fcde",
  1095 => x"c180f750",
  1096 => x"c140e9c3",
  1097 => x"ce78e0dd",
  1098 => x"f8dec187",
  1099 => x"d9ddc148",
  1100 => x"c180fc78",
  1101 => x"2678c8c4",
  1102 => x"5b5e0e4f",
  1103 => x"4c710e5c",
  1104 => x"c192cb4a",
  1105 => x"c882e7dd",
  1106 => x"a2c949a2",
  1107 => x"4b6b974b",
  1108 => x"4969971e",
  1109 => x"1282ca1e",
  1110 => x"e3e8c049",
  1111 => x"d349c087",
  1112 => x"497487f7",
  1113 => x"87eafac0",
  1114 => x"f8f48ef8",
  1115 => x"1e731e87",
  1116 => x"ff494b71",
  1117 => x"497387c3",
  1118 => x"f487fefe",
  1119 => x"731e87e9",
  1120 => x"c64b711e",
  1121 => x"db024aa3",
  1122 => x"028ac187",
  1123 => x"028a87d6",
  1124 => x"8a87dac1",
  1125 => x"87fcc002",
  1126 => x"e1c0028a",
  1127 => x"cb028a87",
  1128 => x"87dbc187",
  1129 => x"c0fd49c7",
  1130 => x"87dec187",
  1131 => x"bfe0ebc2",
  1132 => x"87cbc102",
  1133 => x"c288c148",
  1134 => x"c158e4eb",
  1135 => x"ebc287c1",
  1136 => x"c002bfe4",
  1137 => x"ebc287f9",
  1138 => x"c148bfe0",
  1139 => x"e4ebc280",
  1140 => x"87ebc058",
  1141 => x"bfe0ebc2",
  1142 => x"c289c649",
  1143 => x"c059e4eb",
  1144 => x"da03a9b7",
  1145 => x"e0ebc287",
  1146 => x"d278c048",
  1147 => x"e4ebc287",
  1148 => x"87cb02bf",
  1149 => x"bfe0ebc2",
  1150 => x"c280c648",
  1151 => x"c058e4eb",
  1152 => x"87d5d149",
  1153 => x"f8c04973",
  1154 => x"daf287c8",
  1155 => x"5b5e0e87",
  1156 => x"4c710e5c",
  1157 => x"741e66cc",
  1158 => x"c193cb4b",
  1159 => x"c483e7dd",
  1160 => x"496a4aa3",
  1161 => x"87d0fafe",
  1162 => x"7be7c2c1",
  1163 => x"d449a3c8",
  1164 => x"a3c95166",
  1165 => x"5166d849",
  1166 => x"dc49a3ca",
  1167 => x"f1265166",
  1168 => x"5e0e87e3",
  1169 => x"0e5d5c5b",
  1170 => x"d886d0ff",
  1171 => x"a6c459a6",
  1172 => x"c478c048",
  1173 => x"66c4c180",
  1174 => x"c180c478",
  1175 => x"c180c478",
  1176 => x"e4ebc278",
  1177 => x"c278c148",
  1178 => x"48bfdceb",
  1179 => x"cb05a8de",
  1180 => x"87e5f387",
  1181 => x"a6c84970",
  1182 => x"87e6ce59",
  1183 => x"e987ede8",
  1184 => x"dce887cf",
  1185 => x"c04c7087",
  1186 => x"c102acfb",
  1187 => x"66d487d0",
  1188 => x"87c2c105",
  1189 => x"c11e1ec0",
  1190 => x"dadfc11e",
  1191 => x"fd49c01e",
  1192 => x"d0c187eb",
  1193 => x"82c44a66",
  1194 => x"81c7496a",
  1195 => x"1ec15174",
  1196 => x"496a1ed8",
  1197 => x"ece881c8",
  1198 => x"c186d887",
  1199 => x"c04866c4",
  1200 => x"87c701a8",
  1201 => x"c148a6c4",
  1202 => x"c187ce78",
  1203 => x"c14866c4",
  1204 => x"58a6cc88",
  1205 => x"f8e787c3",
  1206 => x"48a6cc87",
  1207 => x"9c7478c2",
  1208 => x"87facc02",
  1209 => x"c14866c4",
  1210 => x"03a866c8",
  1211 => x"d887efcc",
  1212 => x"78c048a6",
  1213 => x"78c080c4",
  1214 => x"7087e6e6",
  1215 => x"acd0c14c",
  1216 => x"87d7c205",
  1217 => x"e97e66dc",
  1218 => x"497087ca",
  1219 => x"59a6e0c0",
  1220 => x"7087cee6",
  1221 => x"acecc04c",
  1222 => x"87eac105",
  1223 => x"cb4966c4",
  1224 => x"66c0c191",
  1225 => x"4aa1c481",
  1226 => x"a1c84d6a",
  1227 => x"5266dc4a",
  1228 => x"79e9c3c1",
  1229 => x"7087eae5",
  1230 => x"d8029c4c",
  1231 => x"acfbc087",
  1232 => x"7487d202",
  1233 => x"87d9e555",
  1234 => x"029c4c70",
  1235 => x"fbc087c7",
  1236 => x"eeff05ac",
  1237 => x"55e0c087",
  1238 => x"c055c1c2",
  1239 => x"66d47d97",
  1240 => x"05a96e49",
  1241 => x"66c487db",
  1242 => x"a866c848",
  1243 => x"c487ca04",
  1244 => x"80c14866",
  1245 => x"c858a6c8",
  1246 => x"4866c887",
  1247 => x"a6cc88c1",
  1248 => x"87dde458",
  1249 => x"d0c14c70",
  1250 => x"87c805ac",
  1251 => x"c14866d0",
  1252 => x"58a6d480",
  1253 => x"02acd0c1",
  1254 => x"c087e9fd",
  1255 => x"d448a6e0",
  1256 => x"66dc7866",
  1257 => x"66e0c048",
  1258 => x"c3c905a8",
  1259 => x"a6e4c087",
  1260 => x"7e78c048",
  1261 => x"fbc04874",
  1262 => x"a6ecc088",
  1263 => x"02987058",
  1264 => x"4887c8c8",
  1265 => x"ecc088cb",
  1266 => x"987058a6",
  1267 => x"87d0c102",
  1268 => x"c088c948",
  1269 => x"7058a6ec",
  1270 => x"d6c30298",
  1271 => x"88c44887",
  1272 => x"58a6ecc0",
  1273 => x"d0029870",
  1274 => x"88c14887",
  1275 => x"58a6ecc0",
  1276 => x"c2029870",
  1277 => x"ccc787fd",
  1278 => x"48a6d887",
  1279 => x"e278f0c0",
  1280 => x"4c7087df",
  1281 => x"02acecc0",
  1282 => x"dc87c3c0",
  1283 => x"ecc05ca6",
  1284 => x"87cc02ac",
  1285 => x"7087cae2",
  1286 => x"acecc04c",
  1287 => x"87f4ff05",
  1288 => x"02acecc0",
  1289 => x"e187c3c0",
  1290 => x"66d887f7",
  1291 => x"4966d41e",
  1292 => x"4966d41e",
  1293 => x"dadfc11e",
  1294 => x"4966d41e",
  1295 => x"c087cef7",
  1296 => x"dc1eca1e",
  1297 => x"91cb4966",
  1298 => x"8166d8c1",
  1299 => x"c448a6d8",
  1300 => x"66d878a1",
  1301 => x"cce249bf",
  1302 => x"c086d887",
  1303 => x"c106a8b7",
  1304 => x"1ec187c4",
  1305 => x"66c81ede",
  1306 => x"f8e149bf",
  1307 => x"7086c887",
  1308 => x"08c04849",
  1309 => x"58a6dc88",
  1310 => x"06a8b7c0",
  1311 => x"d887e7c0",
  1312 => x"b7dd4866",
  1313 => x"87de03a8",
  1314 => x"d849bf6e",
  1315 => x"e0c08166",
  1316 => x"4966d851",
  1317 => x"bf6e81c1",
  1318 => x"51c1c281",
  1319 => x"c24966d8",
  1320 => x"81bf6e81",
  1321 => x"66cc51c0",
  1322 => x"d080c148",
  1323 => x"7ec158a6",
  1324 => x"e287d8c4",
  1325 => x"a6dc87de",
  1326 => x"87d8e258",
  1327 => x"58a6ecc0",
  1328 => x"05a8ecc0",
  1329 => x"c087cac0",
  1330 => x"d848a6e8",
  1331 => x"c4c07866",
  1332 => x"ccdfff87",
  1333 => x"4966c487",
  1334 => x"c0c191cb",
  1335 => x"80714866",
  1336 => x"4a6e7e70",
  1337 => x"496e82c8",
  1338 => x"66d881ca",
  1339 => x"66e8c051",
  1340 => x"d881c149",
  1341 => x"48c18966",
  1342 => x"49703071",
  1343 => x"977189c1",
  1344 => x"d1efc27a",
  1345 => x"66d849bf",
  1346 => x"4a6a9729",
  1347 => x"c0987148",
  1348 => x"6e58a6f0",
  1349 => x"6981c449",
  1350 => x"66e0c04d",
  1351 => x"a866dc48",
  1352 => x"87c8c002",
  1353 => x"c048a6d8",
  1354 => x"87c5c078",
  1355 => x"c148a6d8",
  1356 => x"1e66d878",
  1357 => x"751ee0c0",
  1358 => x"e8deff49",
  1359 => x"7086c887",
  1360 => x"acb7c04c",
  1361 => x"87d4c106",
  1362 => x"e0c08574",
  1363 => x"75897449",
  1364 => x"d6d9c14b",
  1365 => x"edfe714a",
  1366 => x"85c287ce",
  1367 => x"4866e4c0",
  1368 => x"e8c080c1",
  1369 => x"ecc058a6",
  1370 => x"81c14966",
  1371 => x"c002a970",
  1372 => x"a6d887c8",
  1373 => x"c078c048",
  1374 => x"a6d887c5",
  1375 => x"d878c148",
  1376 => x"a4c21e66",
  1377 => x"48e0c049",
  1378 => x"49708871",
  1379 => x"ff49751e",
  1380 => x"c887d2dd",
  1381 => x"a8b7c086",
  1382 => x"87c0ff01",
  1383 => x"0266e4c0",
  1384 => x"6e87d1c0",
  1385 => x"c081c949",
  1386 => x"6e5166e4",
  1387 => x"f9c4c148",
  1388 => x"87ccc078",
  1389 => x"81c9496e",
  1390 => x"486e51c2",
  1391 => x"78edc5c1",
  1392 => x"c6c07ec1",
  1393 => x"c8dcff87",
  1394 => x"6e4c7087",
  1395 => x"87f5c002",
  1396 => x"c84866c4",
  1397 => x"c004a866",
  1398 => x"66c487cb",
  1399 => x"c880c148",
  1400 => x"e0c058a6",
  1401 => x"4866c887",
  1402 => x"a6cc88c1",
  1403 => x"87d5c058",
  1404 => x"05acc6c1",
  1405 => x"cc87c8c0",
  1406 => x"80c14866",
  1407 => x"ff58a6d0",
  1408 => x"7087cedb",
  1409 => x"4866d04c",
  1410 => x"a6d480c1",
  1411 => x"029c7458",
  1412 => x"c487cbc0",
  1413 => x"c8c14866",
  1414 => x"f304a866",
  1415 => x"daff87d1",
  1416 => x"66c487e6",
  1417 => x"03a8c748",
  1418 => x"c287e5c0",
  1419 => x"c048e4eb",
  1420 => x"4966c478",
  1421 => x"c0c191cb",
  1422 => x"a1c48166",
  1423 => x"c04a6a4a",
  1424 => x"66c47952",
  1425 => x"c880c148",
  1426 => x"a8c758a6",
  1427 => x"87dbff04",
  1428 => x"e18ed0ff",
  1429 => x"203a87cd",
  1430 => x"1e731e00",
  1431 => x"029b4b71",
  1432 => x"ebc287c6",
  1433 => x"78c048e0",
  1434 => x"ebc21ec7",
  1435 => x"1e49bfe0",
  1436 => x"1ee7ddc1",
  1437 => x"bfdcebc2",
  1438 => x"87c6ef49",
  1439 => x"ebc286cc",
  1440 => x"ea49bfdc",
  1441 => x"9b7387cb",
  1442 => x"c187c802",
  1443 => x"c049e7dd",
  1444 => x"e087d1e7",
  1445 => x"731e87d1",
  1446 => x"c24bc01e",
  1447 => x"c048dbdc",
  1448 => x"cadfc150",
  1449 => x"fdc049bf",
  1450 => x"987087c6",
  1451 => x"c187c405",
  1452 => x"734bf9da",
  1453 => x"eedfff48",
  1454 => x"4d4f5287",
  1455 => x"616f6c20",
  1456 => x"676e6964",
  1457 => x"69616620",
  1458 => x"0064656c",
  1459 => x"87e9c71e",
  1460 => x"c4fe49c1",
  1461 => x"e2effe87",
  1462 => x"02987087",
  1463 => x"f8fe87cd",
  1464 => x"987087df",
  1465 => x"c187c402",
  1466 => x"c087c24a",
  1467 => x"059a724a",
  1468 => x"1ec087ce",
  1469 => x"49e0dcc1",
  1470 => x"87edf2c0",
  1471 => x"87fe86c4",
  1472 => x"87c1c1c1",
  1473 => x"dcc11ec0",
  1474 => x"f2c049eb",
  1475 => x"1ec087db",
  1476 => x"7087c3fe",
  1477 => x"d0f2c049",
  1478 => x"87dcc387",
  1479 => x"4f268ef8",
  1480 => x"66204453",
  1481 => x"656c6961",
  1482 => x"42002e64",
  1483 => x"69746f6f",
  1484 => x"2e2e676e",
  1485 => x"c01e002e",
  1486 => x"c087c5e9",
  1487 => x"f687e0f5",
  1488 => x"1e4f2687",
  1489 => x"48e0ebc2",
  1490 => x"ebc278c0",
  1491 => x"78c048dc",
  1492 => x"e187f9fd",
  1493 => x"2648c087",
  1494 => x"4520804f",
  1495 => x"00746978",
  1496 => x"61422080",
  1497 => x"e9006b63",
  1498 => x"f5000010",
  1499 => x"0000002a",
  1500 => x"10e90000",
  1501 => x"2b130000",
  1502 => x"00000000",
  1503 => x"0010e900",
  1504 => x"002b3100",
  1505 => x"00000000",
  1506 => x"000010e9",
  1507 => x"00002b4f",
  1508 => x"e9000000",
  1509 => x"6d000010",
  1510 => x"0000002b",
  1511 => x"10e90000",
  1512 => x"2b8b0000",
  1513 => x"00000000",
  1514 => x"0010e900",
  1515 => x"002ba900",
  1516 => x"00000000",
  1517 => x"000010e9",
  1518 => x"00000000",
  1519 => x"7e000000",
  1520 => x"00000011",
  1521 => x"00000000",
  1522 => x"17ce0000",
  1523 => x"454e0000",
  1524 => x"4f45474f",
  1525 => x"4f522020",
  1526 => x"6f4c004d",
  1527 => x"2a206461",
  1528 => x"fe1e002e",
  1529 => x"78c048f0",
  1530 => x"097909cd",
  1531 => x"1e1e4f26",
  1532 => x"7ebff0fe",
  1533 => x"4f262648",
  1534 => x"48f0fe1e",
  1535 => x"4f2678c1",
  1536 => x"48f0fe1e",
  1537 => x"4f2678c0",
  1538 => x"c04a711e",
  1539 => x"4f265252",
  1540 => x"5c5b5e0e",
  1541 => x"86f40e5d",
  1542 => x"6d974d71",
  1543 => x"4ca5c17e",
  1544 => x"c8486c97",
  1545 => x"486e58a6",
  1546 => x"05a866c4",
  1547 => x"48ff87c5",
  1548 => x"ff87e6c0",
  1549 => x"a5c287ca",
  1550 => x"4b6c9749",
  1551 => x"974ba371",
  1552 => x"6c974b6b",
  1553 => x"c1486e7e",
  1554 => x"58a6c880",
  1555 => x"a6cc98c7",
  1556 => x"7c977058",
  1557 => x"7387e1fe",
  1558 => x"268ef448",
  1559 => x"264c264d",
  1560 => x"0e4f264b",
  1561 => x"0e5c5b5e",
  1562 => x"4c7186f4",
  1563 => x"c34a66d8",
  1564 => x"a4c29aff",
  1565 => x"496c974b",
  1566 => x"7249a173",
  1567 => x"7e6c9751",
  1568 => x"80c1486e",
  1569 => x"c758a6c8",
  1570 => x"58a6cc98",
  1571 => x"8ef45470",
  1572 => x"1e87caff",
  1573 => x"87e8fd1e",
  1574 => x"494abfe0",
  1575 => x"99c0e0c0",
  1576 => x"7287cb02",
  1577 => x"c7efc21e",
  1578 => x"87f7fe49",
  1579 => x"fdfc86c4",
  1580 => x"fd7e7087",
  1581 => x"262687c2",
  1582 => x"efc21e4f",
  1583 => x"c7fd49c7",
  1584 => x"d3e2c187",
  1585 => x"87dafc49",
  1586 => x"2687d5c6",
  1587 => x"5b5e0e4f",
  1588 => x"c20e5d5c",
  1589 => x"4abfe6ef",
  1590 => x"bfe1e4c1",
  1591 => x"bc724c49",
  1592 => x"dbfc4d71",
  1593 => x"744bc087",
  1594 => x"0299d049",
  1595 => x"497587d5",
  1596 => x"1e7199d0",
  1597 => x"ebc11ec0",
  1598 => x"82734aef",
  1599 => x"cac14912",
  1600 => x"c186c887",
  1601 => x"c8832d2c",
  1602 => x"daff04ab",
  1603 => x"87e8fb87",
  1604 => x"48e1e4c1",
  1605 => x"bfe6efc2",
  1606 => x"264d2678",
  1607 => x"264b264c",
  1608 => x"0000004f",
  1609 => x"1e731e00",
  1610 => x"4ac04b71",
  1611 => x"49efebc1",
  1612 => x"69978172",
  1613 => x"05a97349",
  1614 => x"48c187c4",
  1615 => x"82c187ca",
  1616 => x"04aab7c8",
  1617 => x"48c087e6",
  1618 => x"1e87d2ff",
  1619 => x"4b711e73",
  1620 => x"87d1ff49",
  1621 => x"c0029870",
  1622 => x"d0ff87ec",
  1623 => x"78e1c848",
  1624 => x"c548d4ff",
  1625 => x"0266c878",
  1626 => x"e0c387c3",
  1627 => x"0266cc78",
  1628 => x"d4ff87c6",
  1629 => x"78f0c348",
  1630 => x"7348d4ff",
  1631 => x"48d0ff78",
  1632 => x"c078e1c8",
  1633 => x"d4fe78e0",
  1634 => x"5b5e0e87",
  1635 => x"4c710e5c",
  1636 => x"49c7efc2",
  1637 => x"7087f9f9",
  1638 => x"aab7c04a",
  1639 => x"87e3c204",
  1640 => x"05aae0c3",
  1641 => x"e9c187c9",
  1642 => x"78c148cc",
  1643 => x"c387d4c2",
  1644 => x"c905aaf0",
  1645 => x"c8e9c187",
  1646 => x"c178c148",
  1647 => x"e9c187f5",
  1648 => x"c702bfcc",
  1649 => x"c24b7287",
  1650 => x"87c2b3c0",
  1651 => x"9c744b72",
  1652 => x"c187d105",
  1653 => x"1ebfc8e9",
  1654 => x"bfcce9c1",
  1655 => x"fd49721e",
  1656 => x"86c887e9",
  1657 => x"bfc8e9c1",
  1658 => x"87e0c002",
  1659 => x"b7c44973",
  1660 => x"eac19129",
  1661 => x"4a7381ef",
  1662 => x"92c29acf",
  1663 => x"307248c1",
  1664 => x"baff4a70",
  1665 => x"98694872",
  1666 => x"87db7970",
  1667 => x"b7c44973",
  1668 => x"eac19129",
  1669 => x"4a7381ef",
  1670 => x"92c29acf",
  1671 => x"307248c3",
  1672 => x"69484a70",
  1673 => x"c17970b0",
  1674 => x"c048cce9",
  1675 => x"c8e9c178",
  1676 => x"c278c048",
  1677 => x"f749c7ef",
  1678 => x"4a7087d6",
  1679 => x"03aab7c0",
  1680 => x"c087ddfd",
  1681 => x"87d3fb48",
  1682 => x"00000000",
  1683 => x"00000000",
  1684 => x"711e731e",
  1685 => x"87f5f94b",
  1686 => x"ecfc4973",
  1687 => x"87fdfa87",
  1688 => x"724ac01e",
  1689 => x"c191c449",
  1690 => x"c081efea",
  1691 => x"d082c179",
  1692 => x"ee04aab7",
  1693 => x"0e4f2687",
  1694 => x"5d5c5b5e",
  1695 => x"f54d710e",
  1696 => x"4a7587fe",
  1697 => x"922ab7c4",
  1698 => x"82efeac1",
  1699 => x"9ccf4c75",
  1700 => x"496a94c2",
  1701 => x"c32b744b",
  1702 => x"7448c29b",
  1703 => x"ff4c7030",
  1704 => x"714874bc",
  1705 => x"f57a7098",
  1706 => x"487387ce",
  1707 => x"0087eaf9",
  1708 => x"00000000",
  1709 => x"00000000",
  1710 => x"00000000",
  1711 => x"00000000",
  1712 => x"00000000",
  1713 => x"00000000",
  1714 => x"00000000",
  1715 => x"00000000",
  1716 => x"00000000",
  1717 => x"00000000",
  1718 => x"00000000",
  1719 => x"00000000",
  1720 => x"00000000",
  1721 => x"00000000",
  1722 => x"00000000",
  1723 => x"16000000",
  1724 => x"2e25261e",
  1725 => x"1e3e3d36",
  1726 => x"c848d0ff",
  1727 => x"487178e1",
  1728 => x"7808d4ff",
  1729 => x"ff1e4f26",
  1730 => x"e1c848d0",
  1731 => x"ff487178",
  1732 => x"c47808d4",
  1733 => x"d4ff4866",
  1734 => x"4f267808",
  1735 => x"c44a711e",
  1736 => x"721e4966",
  1737 => x"87deff49",
  1738 => x"c048d0ff",
  1739 => x"262678e0",
  1740 => x"4a711e4f",
  1741 => x"c11e66c4",
  1742 => x"ff49a2e0",
  1743 => x"66c887c8",
  1744 => x"29b7c849",
  1745 => x"7148d4ff",
  1746 => x"48d0ff78",
  1747 => x"2678e0c0",
  1748 => x"ff1e4f26",
  1749 => x"ffc34ad4",
  1750 => x"48d0ff7a",
  1751 => x"de78e1c8",
  1752 => x"d1efc27a",
  1753 => x"48497abf",
  1754 => x"7a7028c8",
  1755 => x"28d04871",
  1756 => x"48717a70",
  1757 => x"7a7028d8",
  1758 => x"c048d0ff",
  1759 => x"4f2678e0",
  1760 => x"5c5b5e0e",
  1761 => x"4c710e5d",
  1762 => x"bfd1efc2",
  1763 => x"2b744b4d",
  1764 => x"c19b66d0",
  1765 => x"ab66d483",
  1766 => x"c087c204",
  1767 => x"d04a744b",
  1768 => x"31724966",
  1769 => x"9975b9ff",
  1770 => x"30724873",
  1771 => x"71484a70",
  1772 => x"d5efc2b0",
  1773 => x"87dafe58",
  1774 => x"4c264d26",
  1775 => x"4f264b26",
  1776 => x"48d0ff1e",
  1777 => x"7178c9c8",
  1778 => x"08d4ff48",
  1779 => x"1e4f2678",
  1780 => x"eb494a71",
  1781 => x"48d0ff87",
  1782 => x"4f2678c8",
  1783 => x"711e731e",
  1784 => x"e1efc24b",
  1785 => x"87c302bf",
  1786 => x"ff87ebc2",
  1787 => x"c9c848d0",
  1788 => x"c0497378",
  1789 => x"d4ffb1e0",
  1790 => x"c2787148",
  1791 => x"c048d5ef",
  1792 => x"0266c878",
  1793 => x"ffc387c5",
  1794 => x"c087c249",
  1795 => x"ddefc249",
  1796 => x"0266cc59",
  1797 => x"d5c587c6",
  1798 => x"87c44ad5",
  1799 => x"4affffcf",
  1800 => x"5ae1efc2",
  1801 => x"48e1efc2",
  1802 => x"87c478c1",
  1803 => x"4c264d26",
  1804 => x"4f264b26",
  1805 => x"5c5b5e0e",
  1806 => x"4a710e5d",
  1807 => x"bfddefc2",
  1808 => x"029a724c",
  1809 => x"c84987cb",
  1810 => x"d2efc191",
  1811 => x"c483714b",
  1812 => x"d2f3c187",
  1813 => x"134dc04b",
  1814 => x"c2997449",
  1815 => x"b9bfd9ef",
  1816 => x"7148d4ff",
  1817 => x"2cb7c178",
  1818 => x"adb7c885",
  1819 => x"c287e804",
  1820 => x"48bfd5ef",
  1821 => x"efc280c8",
  1822 => x"effe58d9",
  1823 => x"1e731e87",
  1824 => x"4a134b71",
  1825 => x"87cb029a",
  1826 => x"e7fe4972",
  1827 => x"9a4a1387",
  1828 => x"fe87f505",
  1829 => x"c21e87da",
  1830 => x"49bfd5ef",
  1831 => x"48d5efc2",
  1832 => x"c478a1c1",
  1833 => x"03a9b7c0",
  1834 => x"d4ff87db",
  1835 => x"d9efc248",
  1836 => x"efc278bf",
  1837 => x"c249bfd5",
  1838 => x"c148d5ef",
  1839 => x"c0c478a1",
  1840 => x"e504a9b7",
  1841 => x"48d0ff87",
  1842 => x"efc278c8",
  1843 => x"78c048e1",
  1844 => x"00004f26",
  1845 => x"00000000",
  1846 => x"00000000",
  1847 => x"005f5f00",
  1848 => x"03000000",
  1849 => x"03030003",
  1850 => x"7f140000",
  1851 => x"7f7f147f",
  1852 => x"24000014",
  1853 => x"3a6b6b2e",
  1854 => x"6a4c0012",
  1855 => x"566c1836",
  1856 => x"7e300032",
  1857 => x"3a77594f",
  1858 => x"00004068",
  1859 => x"00030704",
  1860 => x"00000000",
  1861 => x"41633e1c",
  1862 => x"00000000",
  1863 => x"1c3e6341",
  1864 => x"2a080000",
  1865 => x"3e1c1c3e",
  1866 => x"0800082a",
  1867 => x"083e3e08",
  1868 => x"00000008",
  1869 => x"0060e080",
  1870 => x"08000000",
  1871 => x"08080808",
  1872 => x"00000008",
  1873 => x"00606000",
  1874 => x"60400000",
  1875 => x"060c1830",
  1876 => x"3e000103",
  1877 => x"7f4d597f",
  1878 => x"0400003e",
  1879 => x"007f7f06",
  1880 => x"42000000",
  1881 => x"4f597163",
  1882 => x"22000046",
  1883 => x"7f494963",
  1884 => x"1c180036",
  1885 => x"7f7f1316",
  1886 => x"27000010",
  1887 => x"7d454567",
  1888 => x"3c000039",
  1889 => x"79494b7e",
  1890 => x"01000030",
  1891 => x"0f797101",
  1892 => x"36000007",
  1893 => x"7f49497f",
  1894 => x"06000036",
  1895 => x"3f69494f",
  1896 => x"0000001e",
  1897 => x"00666600",
  1898 => x"00000000",
  1899 => x"0066e680",
  1900 => x"08000000",
  1901 => x"22141408",
  1902 => x"14000022",
  1903 => x"14141414",
  1904 => x"22000014",
  1905 => x"08141422",
  1906 => x"02000008",
  1907 => x"0f595103",
  1908 => x"7f3e0006",
  1909 => x"1f555d41",
  1910 => x"7e00001e",
  1911 => x"7f09097f",
  1912 => x"7f00007e",
  1913 => x"7f49497f",
  1914 => x"1c000036",
  1915 => x"4141633e",
  1916 => x"7f000041",
  1917 => x"3e63417f",
  1918 => x"7f00001c",
  1919 => x"4149497f",
  1920 => x"7f000041",
  1921 => x"0109097f",
  1922 => x"3e000001",
  1923 => x"7b49417f",
  1924 => x"7f00007a",
  1925 => x"7f08087f",
  1926 => x"0000007f",
  1927 => x"417f7f41",
  1928 => x"20000000",
  1929 => x"7f404060",
  1930 => x"7f7f003f",
  1931 => x"63361c08",
  1932 => x"7f000041",
  1933 => x"4040407f",
  1934 => x"7f7f0040",
  1935 => x"7f060c06",
  1936 => x"7f7f007f",
  1937 => x"7f180c06",
  1938 => x"3e00007f",
  1939 => x"7f41417f",
  1940 => x"7f00003e",
  1941 => x"0f09097f",
  1942 => x"7f3e0006",
  1943 => x"7e7f6141",
  1944 => x"7f000040",
  1945 => x"7f19097f",
  1946 => x"26000066",
  1947 => x"7b594d6f",
  1948 => x"01000032",
  1949 => x"017f7f01",
  1950 => x"3f000001",
  1951 => x"7f40407f",
  1952 => x"0f00003f",
  1953 => x"3f70703f",
  1954 => x"7f7f000f",
  1955 => x"7f301830",
  1956 => x"6341007f",
  1957 => x"361c1c36",
  1958 => x"03014163",
  1959 => x"067c7c06",
  1960 => x"71610103",
  1961 => x"43474d59",
  1962 => x"00000041",
  1963 => x"41417f7f",
  1964 => x"03010000",
  1965 => x"30180c06",
  1966 => x"00004060",
  1967 => x"7f7f4141",
  1968 => x"0c080000",
  1969 => x"0c060306",
  1970 => x"80800008",
  1971 => x"80808080",
  1972 => x"00000080",
  1973 => x"04070300",
  1974 => x"20000000",
  1975 => x"7c545474",
  1976 => x"7f000078",
  1977 => x"7c44447f",
  1978 => x"38000038",
  1979 => x"4444447c",
  1980 => x"38000000",
  1981 => x"7f44447c",
  1982 => x"3800007f",
  1983 => x"5c54547c",
  1984 => x"04000018",
  1985 => x"05057f7e",
  1986 => x"18000000",
  1987 => x"fca4a4bc",
  1988 => x"7f00007c",
  1989 => x"7c04047f",
  1990 => x"00000078",
  1991 => x"407d3d00",
  1992 => x"80000000",
  1993 => x"7dfd8080",
  1994 => x"7f000000",
  1995 => x"6c38107f",
  1996 => x"00000044",
  1997 => x"407f3f00",
  1998 => x"7c7c0000",
  1999 => x"7c0c180c",
  2000 => x"7c000078",
  2001 => x"7c04047c",
  2002 => x"38000078",
  2003 => x"7c44447c",
  2004 => x"fc000038",
  2005 => x"3c2424fc",
  2006 => x"18000018",
  2007 => x"fc24243c",
  2008 => x"7c0000fc",
  2009 => x"0c04047c",
  2010 => x"48000008",
  2011 => x"7454545c",
  2012 => x"04000020",
  2013 => x"44447f3f",
  2014 => x"3c000000",
  2015 => x"7c40407c",
  2016 => x"1c00007c",
  2017 => x"3c60603c",
  2018 => x"7c3c001c",
  2019 => x"7c603060",
  2020 => x"6c44003c",
  2021 => x"6c381038",
  2022 => x"1c000044",
  2023 => x"3c60e0bc",
  2024 => x"4400001c",
  2025 => x"4c5c7464",
  2026 => x"08000044",
  2027 => x"41773e08",
  2028 => x"00000041",
  2029 => x"007f7f00",
  2030 => x"41000000",
  2031 => x"083e7741",
  2032 => x"01020008",
  2033 => x"02020301",
  2034 => x"7f7f0001",
  2035 => x"7f7f7f7f",
  2036 => x"0808007f",
  2037 => x"3e3e1c1c",
  2038 => x"7f7f7f7f",
  2039 => x"1c1c3e3e",
  2040 => x"10000808",
  2041 => x"187c7c18",
  2042 => x"10000010",
  2043 => x"307c7c30",
  2044 => x"30100010",
  2045 => x"1e786060",
  2046 => x"66420006",
  2047 => x"663c183c",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
