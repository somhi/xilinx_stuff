
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"e4",x"f0",x"c2",x"87"),
    12 => (x"86",x"c0",x"c6",x"4e"),
    13 => (x"49",x"e4",x"f0",x"c2"),
    14 => (x"48",x"c4",x"de",x"c2"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"f8",x"db"),
    19 => (x"1e",x"87",x"fc",x"98"),
    20 => (x"1e",x"73",x"1e",x"72"),
    21 => (x"02",x"11",x"48",x"12"),
    22 => (x"c3",x"4b",x"87",x"ca"),
    23 => (x"73",x"9b",x"98",x"df"),
    24 => (x"87",x"f0",x"02",x"88"),
    25 => (x"4a",x"26",x"4b",x"26"),
    26 => (x"73",x"1e",x"4f",x"26"),
    27 => (x"c1",x"1e",x"72",x"1e"),
    28 => (x"87",x"ca",x"04",x"8b"),
    29 => (x"02",x"11",x"48",x"12"),
    30 => (x"02",x"88",x"87",x"c4"),
    31 => (x"4a",x"26",x"87",x"f1"),
    32 => (x"4f",x"26",x"4b",x"26"),
    33 => (x"73",x"1e",x"74",x"1e"),
    34 => (x"c1",x"1e",x"72",x"1e"),
    35 => (x"87",x"d0",x"04",x"8b"),
    36 => (x"02",x"11",x"48",x"12"),
    37 => (x"c3",x"4c",x"87",x"ca"),
    38 => (x"74",x"9c",x"98",x"df"),
    39 => (x"87",x"eb",x"02",x"88"),
    40 => (x"4b",x"26",x"4a",x"26"),
    41 => (x"4f",x"26",x"4c",x"26"),
    42 => (x"81",x"48",x"73",x"1e"),
    43 => (x"c5",x"02",x"a9",x"73"),
    44 => (x"05",x"53",x"12",x"87"),
    45 => (x"4f",x"26",x"87",x"f6"),
    46 => (x"4a",x"66",x"c4",x"1e"),
    47 => (x"51",x"12",x"48",x"71"),
    48 => (x"26",x"87",x"fb",x"05"),
    49 => (x"48",x"11",x"1e",x"4f"),
    50 => (x"78",x"08",x"d4",x"ff"),
    51 => (x"c1",x"48",x"66",x"c4"),
    52 => (x"58",x"a6",x"c8",x"88"),
    53 => (x"ed",x"05",x"98",x"70"),
    54 => (x"1e",x"4f",x"26",x"87"),
    55 => (x"c3",x"48",x"d4",x"ff"),
    56 => (x"51",x"68",x"78",x"ff"),
    57 => (x"c1",x"48",x"66",x"c4"),
    58 => (x"58",x"a6",x"c8",x"88"),
    59 => (x"eb",x"05",x"98",x"70"),
    60 => (x"1e",x"4f",x"26",x"87"),
    61 => (x"d4",x"ff",x"1e",x"73"),
    62 => (x"7b",x"ff",x"c3",x"4b"),
    63 => (x"ff",x"c3",x"4a",x"6b"),
    64 => (x"c8",x"49",x"6b",x"7b"),
    65 => (x"c3",x"b1",x"72",x"32"),
    66 => (x"4a",x"6b",x"7b",x"ff"),
    67 => (x"b2",x"71",x"31",x"c8"),
    68 => (x"6b",x"7b",x"ff",x"c3"),
    69 => (x"72",x"32",x"c8",x"49"),
    70 => (x"c4",x"48",x"71",x"b1"),
    71 => (x"26",x"4d",x"26",x"87"),
    72 => (x"26",x"4b",x"26",x"4c"),
    73 => (x"5b",x"5e",x"0e",x"4f"),
    74 => (x"71",x"0e",x"5d",x"5c"),
    75 => (x"4c",x"d4",x"ff",x"4a"),
    76 => (x"ff",x"c3",x"49",x"72"),
    77 => (x"c2",x"7c",x"71",x"99"),
    78 => (x"05",x"bf",x"c4",x"de"),
    79 => (x"66",x"d0",x"87",x"c8"),
    80 => (x"d4",x"30",x"c9",x"48"),
    81 => (x"66",x"d0",x"58",x"a6"),
    82 => (x"c3",x"29",x"d8",x"49"),
    83 => (x"7c",x"71",x"99",x"ff"),
    84 => (x"d0",x"49",x"66",x"d0"),
    85 => (x"99",x"ff",x"c3",x"29"),
    86 => (x"66",x"d0",x"7c",x"71"),
    87 => (x"c3",x"29",x"c8",x"49"),
    88 => (x"7c",x"71",x"99",x"ff"),
    89 => (x"c3",x"49",x"66",x"d0"),
    90 => (x"7c",x"71",x"99",x"ff"),
    91 => (x"29",x"d0",x"49",x"72"),
    92 => (x"71",x"99",x"ff",x"c3"),
    93 => (x"c9",x"4b",x"6c",x"7c"),
    94 => (x"c3",x"4d",x"ff",x"f0"),
    95 => (x"d0",x"05",x"ab",x"ff"),
    96 => (x"7c",x"ff",x"c3",x"87"),
    97 => (x"8d",x"c1",x"4b",x"6c"),
    98 => (x"c3",x"87",x"c6",x"02"),
    99 => (x"f0",x"02",x"ab",x"ff"),
   100 => (x"fe",x"48",x"73",x"87"),
   101 => (x"c0",x"1e",x"87",x"c7"),
   102 => (x"48",x"d4",x"ff",x"49"),
   103 => (x"c1",x"78",x"ff",x"c3"),
   104 => (x"b7",x"c8",x"c3",x"81"),
   105 => (x"87",x"f1",x"04",x"a9"),
   106 => (x"73",x"1e",x"4f",x"26"),
   107 => (x"c4",x"87",x"e7",x"1e"),
   108 => (x"c0",x"4b",x"df",x"f8"),
   109 => (x"f0",x"ff",x"c0",x"1e"),
   110 => (x"fd",x"49",x"f7",x"c1"),
   111 => (x"86",x"c4",x"87",x"e7"),
   112 => (x"c0",x"05",x"a8",x"c1"),
   113 => (x"d4",x"ff",x"87",x"ea"),
   114 => (x"78",x"ff",x"c3",x"48"),
   115 => (x"c0",x"c0",x"c0",x"c1"),
   116 => (x"c0",x"1e",x"c0",x"c0"),
   117 => (x"e9",x"c1",x"f0",x"e1"),
   118 => (x"87",x"c9",x"fd",x"49"),
   119 => (x"98",x"70",x"86",x"c4"),
   120 => (x"ff",x"87",x"ca",x"05"),
   121 => (x"ff",x"c3",x"48",x"d4"),
   122 => (x"cb",x"48",x"c1",x"78"),
   123 => (x"87",x"e6",x"fe",x"87"),
   124 => (x"fe",x"05",x"8b",x"c1"),
   125 => (x"48",x"c0",x"87",x"fd"),
   126 => (x"1e",x"87",x"e6",x"fc"),
   127 => (x"d4",x"ff",x"1e",x"73"),
   128 => (x"78",x"ff",x"c3",x"48"),
   129 => (x"1e",x"c0",x"4b",x"d3"),
   130 => (x"c1",x"f0",x"ff",x"c0"),
   131 => (x"d4",x"fc",x"49",x"c1"),
   132 => (x"70",x"86",x"c4",x"87"),
   133 => (x"87",x"ca",x"05",x"98"),
   134 => (x"c3",x"48",x"d4",x"ff"),
   135 => (x"48",x"c1",x"78",x"ff"),
   136 => (x"f1",x"fd",x"87",x"cb"),
   137 => (x"05",x"8b",x"c1",x"87"),
   138 => (x"c0",x"87",x"db",x"ff"),
   139 => (x"87",x"f1",x"fb",x"48"),
   140 => (x"5c",x"5b",x"5e",x"0e"),
   141 => (x"4c",x"d4",x"ff",x"0e"),
   142 => (x"c6",x"87",x"db",x"fd"),
   143 => (x"e1",x"c0",x"1e",x"ea"),
   144 => (x"49",x"c8",x"c1",x"f0"),
   145 => (x"c4",x"87",x"de",x"fb"),
   146 => (x"02",x"a8",x"c1",x"86"),
   147 => (x"ea",x"fe",x"87",x"c8"),
   148 => (x"c1",x"48",x"c0",x"87"),
   149 => (x"da",x"fa",x"87",x"e2"),
   150 => (x"cf",x"49",x"70",x"87"),
   151 => (x"c6",x"99",x"ff",x"ff"),
   152 => (x"c8",x"02",x"a9",x"ea"),
   153 => (x"87",x"d3",x"fe",x"87"),
   154 => (x"cb",x"c1",x"48",x"c0"),
   155 => (x"7c",x"ff",x"c3",x"87"),
   156 => (x"fc",x"4b",x"f1",x"c0"),
   157 => (x"98",x"70",x"87",x"f4"),
   158 => (x"87",x"eb",x"c0",x"02"),
   159 => (x"ff",x"c0",x"1e",x"c0"),
   160 => (x"49",x"fa",x"c1",x"f0"),
   161 => (x"c4",x"87",x"de",x"fa"),
   162 => (x"05",x"98",x"70",x"86"),
   163 => (x"ff",x"c3",x"87",x"d9"),
   164 => (x"c3",x"49",x"6c",x"7c"),
   165 => (x"7c",x"7c",x"7c",x"ff"),
   166 => (x"99",x"c0",x"c1",x"7c"),
   167 => (x"c1",x"87",x"c4",x"02"),
   168 => (x"c0",x"87",x"d5",x"48"),
   169 => (x"c2",x"87",x"d1",x"48"),
   170 => (x"87",x"c4",x"05",x"ab"),
   171 => (x"87",x"c8",x"48",x"c0"),
   172 => (x"fe",x"05",x"8b",x"c1"),
   173 => (x"48",x"c0",x"87",x"fd"),
   174 => (x"1e",x"87",x"e4",x"f9"),
   175 => (x"de",x"c2",x"1e",x"73"),
   176 => (x"78",x"c1",x"48",x"c4"),
   177 => (x"d0",x"ff",x"4b",x"c7"),
   178 => (x"fb",x"78",x"c2",x"48"),
   179 => (x"d0",x"ff",x"87",x"c8"),
   180 => (x"c0",x"78",x"c3",x"48"),
   181 => (x"d0",x"e5",x"c0",x"1e"),
   182 => (x"f9",x"49",x"c0",x"c1"),
   183 => (x"86",x"c4",x"87",x"c7"),
   184 => (x"c1",x"05",x"a8",x"c1"),
   185 => (x"ab",x"c2",x"4b",x"87"),
   186 => (x"c0",x"87",x"c5",x"05"),
   187 => (x"87",x"f9",x"c0",x"48"),
   188 => (x"ff",x"05",x"8b",x"c1"),
   189 => (x"f7",x"fc",x"87",x"d0"),
   190 => (x"c8",x"de",x"c2",x"87"),
   191 => (x"05",x"98",x"70",x"58"),
   192 => (x"1e",x"c1",x"87",x"cd"),
   193 => (x"c1",x"f0",x"ff",x"c0"),
   194 => (x"d8",x"f8",x"49",x"d0"),
   195 => (x"ff",x"86",x"c4",x"87"),
   196 => (x"ff",x"c3",x"48",x"d4"),
   197 => (x"87",x"e0",x"c4",x"78"),
   198 => (x"58",x"cc",x"de",x"c2"),
   199 => (x"c2",x"48",x"d0",x"ff"),
   200 => (x"48",x"d4",x"ff",x"78"),
   201 => (x"c1",x"78",x"ff",x"c3"),
   202 => (x"87",x"f5",x"f7",x"48"),
   203 => (x"5c",x"5b",x"5e",x"0e"),
   204 => (x"4a",x"71",x"0e",x"5d"),
   205 => (x"ff",x"4d",x"ff",x"c3"),
   206 => (x"7c",x"75",x"4c",x"d4"),
   207 => (x"c4",x"48",x"d0",x"ff"),
   208 => (x"7c",x"75",x"78",x"c3"),
   209 => (x"ff",x"c0",x"1e",x"72"),
   210 => (x"49",x"d8",x"c1",x"f0"),
   211 => (x"c4",x"87",x"d6",x"f7"),
   212 => (x"02",x"98",x"70",x"86"),
   213 => (x"48",x"c0",x"87",x"c5"),
   214 => (x"75",x"87",x"f0",x"c0"),
   215 => (x"7c",x"fe",x"c3",x"7c"),
   216 => (x"d4",x"1e",x"c0",x"c8"),
   217 => (x"dc",x"f5",x"49",x"66"),
   218 => (x"75",x"86",x"c4",x"87"),
   219 => (x"75",x"7c",x"75",x"7c"),
   220 => (x"e0",x"da",x"d8",x"7c"),
   221 => (x"6c",x"7c",x"75",x"4b"),
   222 => (x"c5",x"05",x"99",x"49"),
   223 => (x"05",x"8b",x"c1",x"87"),
   224 => (x"7c",x"75",x"87",x"f3"),
   225 => (x"c2",x"48",x"d0",x"ff"),
   226 => (x"f6",x"48",x"c1",x"78"),
   227 => (x"ff",x"1e",x"87",x"cf"),
   228 => (x"d0",x"ff",x"4a",x"d4"),
   229 => (x"78",x"d1",x"c4",x"48"),
   230 => (x"c1",x"7a",x"ff",x"c3"),
   231 => (x"87",x"f8",x"05",x"89"),
   232 => (x"73",x"1e",x"4f",x"26"),
   233 => (x"c5",x"4b",x"71",x"1e"),
   234 => (x"4a",x"df",x"cd",x"ee"),
   235 => (x"c3",x"48",x"d4",x"ff"),
   236 => (x"48",x"68",x"78",x"ff"),
   237 => (x"02",x"a8",x"fe",x"c3"),
   238 => (x"8a",x"c1",x"87",x"c5"),
   239 => (x"72",x"87",x"ed",x"05"),
   240 => (x"87",x"c5",x"05",x"9a"),
   241 => (x"ea",x"c0",x"48",x"c0"),
   242 => (x"02",x"9b",x"73",x"87"),
   243 => (x"66",x"c8",x"87",x"cc"),
   244 => (x"f4",x"49",x"73",x"1e"),
   245 => (x"86",x"c4",x"87",x"c5"),
   246 => (x"66",x"c8",x"87",x"c6"),
   247 => (x"87",x"ee",x"fe",x"49"),
   248 => (x"c3",x"48",x"d4",x"ff"),
   249 => (x"73",x"78",x"78",x"ff"),
   250 => (x"87",x"c5",x"05",x"9b"),
   251 => (x"d0",x"48",x"d0",x"ff"),
   252 => (x"f4",x"48",x"c1",x"78"),
   253 => (x"73",x"1e",x"87",x"eb"),
   254 => (x"c0",x"4a",x"71",x"1e"),
   255 => (x"48",x"d4",x"ff",x"4b"),
   256 => (x"ff",x"78",x"ff",x"c3"),
   257 => (x"c3",x"c4",x"48",x"d0"),
   258 => (x"48",x"d4",x"ff",x"78"),
   259 => (x"72",x"78",x"ff",x"c3"),
   260 => (x"f0",x"ff",x"c0",x"1e"),
   261 => (x"f4",x"49",x"d1",x"c1"),
   262 => (x"86",x"c4",x"87",x"cb"),
   263 => (x"cd",x"05",x"98",x"70"),
   264 => (x"1e",x"c0",x"c8",x"87"),
   265 => (x"fd",x"49",x"66",x"cc"),
   266 => (x"86",x"c4",x"87",x"f8"),
   267 => (x"d0",x"ff",x"4b",x"70"),
   268 => (x"73",x"78",x"c2",x"48"),
   269 => (x"87",x"e9",x"f3",x"48"),
   270 => (x"5c",x"5b",x"5e",x"0e"),
   271 => (x"1e",x"c0",x"0e",x"5d"),
   272 => (x"c1",x"f0",x"ff",x"c0"),
   273 => (x"dc",x"f3",x"49",x"c9"),
   274 => (x"c2",x"1e",x"d2",x"87"),
   275 => (x"fd",x"49",x"cc",x"de"),
   276 => (x"86",x"c8",x"87",x"d0"),
   277 => (x"84",x"c1",x"4c",x"c0"),
   278 => (x"04",x"ac",x"b7",x"d2"),
   279 => (x"de",x"c2",x"87",x"f8"),
   280 => (x"49",x"bf",x"97",x"cc"),
   281 => (x"c1",x"99",x"c0",x"c3"),
   282 => (x"c0",x"05",x"a9",x"c0"),
   283 => (x"de",x"c2",x"87",x"e7"),
   284 => (x"49",x"bf",x"97",x"d3"),
   285 => (x"de",x"c2",x"31",x"d0"),
   286 => (x"4a",x"bf",x"97",x"d4"),
   287 => (x"b1",x"72",x"32",x"c8"),
   288 => (x"97",x"d5",x"de",x"c2"),
   289 => (x"71",x"b1",x"4a",x"bf"),
   290 => (x"ff",x"ff",x"cf",x"4c"),
   291 => (x"84",x"c1",x"9c",x"ff"),
   292 => (x"e7",x"c1",x"34",x"ca"),
   293 => (x"d5",x"de",x"c2",x"87"),
   294 => (x"c1",x"49",x"bf",x"97"),
   295 => (x"c2",x"99",x"c6",x"31"),
   296 => (x"bf",x"97",x"d6",x"de"),
   297 => (x"2a",x"b7",x"c7",x"4a"),
   298 => (x"de",x"c2",x"b1",x"72"),
   299 => (x"4a",x"bf",x"97",x"d1"),
   300 => (x"c2",x"9d",x"cf",x"4d"),
   301 => (x"bf",x"97",x"d2",x"de"),
   302 => (x"ca",x"9a",x"c3",x"4a"),
   303 => (x"d3",x"de",x"c2",x"32"),
   304 => (x"c2",x"4b",x"bf",x"97"),
   305 => (x"c2",x"b2",x"73",x"33"),
   306 => (x"bf",x"97",x"d4",x"de"),
   307 => (x"9b",x"c0",x"c3",x"4b"),
   308 => (x"73",x"2b",x"b7",x"c6"),
   309 => (x"c1",x"81",x"c2",x"b2"),
   310 => (x"70",x"30",x"71",x"48"),
   311 => (x"75",x"48",x"c1",x"49"),
   312 => (x"72",x"4d",x"70",x"30"),
   313 => (x"71",x"84",x"c1",x"4c"),
   314 => (x"b7",x"c0",x"c8",x"94"),
   315 => (x"87",x"cc",x"06",x"ad"),
   316 => (x"2d",x"b7",x"34",x"c1"),
   317 => (x"ad",x"b7",x"c0",x"c8"),
   318 => (x"87",x"f4",x"ff",x"01"),
   319 => (x"dc",x"f0",x"48",x"74"),
   320 => (x"5b",x"5e",x"0e",x"87"),
   321 => (x"f8",x"0e",x"5d",x"5c"),
   322 => (x"f2",x"e6",x"c2",x"86"),
   323 => (x"c2",x"78",x"c0",x"48"),
   324 => (x"c0",x"1e",x"ea",x"de"),
   325 => (x"87",x"de",x"fb",x"49"),
   326 => (x"98",x"70",x"86",x"c4"),
   327 => (x"c0",x"87",x"c5",x"05"),
   328 => (x"87",x"ce",x"c9",x"48"),
   329 => (x"7e",x"c1",x"4d",x"c0"),
   330 => (x"bf",x"cb",x"f2",x"c0"),
   331 => (x"e0",x"df",x"c2",x"49"),
   332 => (x"4b",x"c8",x"71",x"4a"),
   333 => (x"70",x"87",x"f3",x"ec"),
   334 => (x"87",x"c2",x"05",x"98"),
   335 => (x"f2",x"c0",x"7e",x"c0"),
   336 => (x"c2",x"49",x"bf",x"c7"),
   337 => (x"71",x"4a",x"fc",x"df"),
   338 => (x"dd",x"ec",x"4b",x"c8"),
   339 => (x"05",x"98",x"70",x"87"),
   340 => (x"7e",x"c0",x"87",x"c2"),
   341 => (x"fd",x"c0",x"02",x"6e"),
   342 => (x"f0",x"e5",x"c2",x"87"),
   343 => (x"e6",x"c2",x"4d",x"bf"),
   344 => (x"7e",x"bf",x"9f",x"e8"),
   345 => (x"ea",x"d6",x"c5",x"48"),
   346 => (x"87",x"c7",x"05",x"a8"),
   347 => (x"bf",x"f0",x"e5",x"c2"),
   348 => (x"6e",x"87",x"ce",x"4d"),
   349 => (x"d5",x"e9",x"ca",x"48"),
   350 => (x"87",x"c5",x"02",x"a8"),
   351 => (x"f1",x"c7",x"48",x"c0"),
   352 => (x"ea",x"de",x"c2",x"87"),
   353 => (x"f9",x"49",x"75",x"1e"),
   354 => (x"86",x"c4",x"87",x"ec"),
   355 => (x"c5",x"05",x"98",x"70"),
   356 => (x"c7",x"48",x"c0",x"87"),
   357 => (x"f2",x"c0",x"87",x"dc"),
   358 => (x"c2",x"49",x"bf",x"c7"),
   359 => (x"71",x"4a",x"fc",x"df"),
   360 => (x"c5",x"eb",x"4b",x"c8"),
   361 => (x"05",x"98",x"70",x"87"),
   362 => (x"e6",x"c2",x"87",x"c8"),
   363 => (x"78",x"c1",x"48",x"f2"),
   364 => (x"f2",x"c0",x"87",x"da"),
   365 => (x"c2",x"49",x"bf",x"cb"),
   366 => (x"71",x"4a",x"e0",x"df"),
   367 => (x"e9",x"ea",x"4b",x"c8"),
   368 => (x"02",x"98",x"70",x"87"),
   369 => (x"c0",x"87",x"c5",x"c0"),
   370 => (x"87",x"e6",x"c6",x"48"),
   371 => (x"97",x"e8",x"e6",x"c2"),
   372 => (x"d5",x"c1",x"49",x"bf"),
   373 => (x"cd",x"c0",x"05",x"a9"),
   374 => (x"e9",x"e6",x"c2",x"87"),
   375 => (x"c2",x"49",x"bf",x"97"),
   376 => (x"c0",x"02",x"a9",x"ea"),
   377 => (x"48",x"c0",x"87",x"c5"),
   378 => (x"c2",x"87",x"c7",x"c6"),
   379 => (x"bf",x"97",x"ea",x"de"),
   380 => (x"e9",x"c3",x"48",x"7e"),
   381 => (x"ce",x"c0",x"02",x"a8"),
   382 => (x"c3",x"48",x"6e",x"87"),
   383 => (x"c0",x"02",x"a8",x"eb"),
   384 => (x"48",x"c0",x"87",x"c5"),
   385 => (x"c2",x"87",x"eb",x"c5"),
   386 => (x"bf",x"97",x"f5",x"de"),
   387 => (x"c0",x"05",x"99",x"49"),
   388 => (x"de",x"c2",x"87",x"cc"),
   389 => (x"49",x"bf",x"97",x"f6"),
   390 => (x"c0",x"02",x"a9",x"c2"),
   391 => (x"48",x"c0",x"87",x"c5"),
   392 => (x"c2",x"87",x"cf",x"c5"),
   393 => (x"bf",x"97",x"f7",x"de"),
   394 => (x"ee",x"e6",x"c2",x"48"),
   395 => (x"48",x"4c",x"70",x"58"),
   396 => (x"e6",x"c2",x"88",x"c1"),
   397 => (x"de",x"c2",x"58",x"f2"),
   398 => (x"49",x"bf",x"97",x"f8"),
   399 => (x"de",x"c2",x"81",x"75"),
   400 => (x"4a",x"bf",x"97",x"f9"),
   401 => (x"a1",x"72",x"32",x"c8"),
   402 => (x"ff",x"ea",x"c2",x"7e"),
   403 => (x"c2",x"78",x"6e",x"48"),
   404 => (x"bf",x"97",x"fa",x"de"),
   405 => (x"58",x"a6",x"c8",x"48"),
   406 => (x"bf",x"f2",x"e6",x"c2"),
   407 => (x"87",x"d4",x"c2",x"02"),
   408 => (x"bf",x"c7",x"f2",x"c0"),
   409 => (x"fc",x"df",x"c2",x"49"),
   410 => (x"4b",x"c8",x"71",x"4a"),
   411 => (x"70",x"87",x"fb",x"e7"),
   412 => (x"c5",x"c0",x"02",x"98"),
   413 => (x"c3",x"48",x"c0",x"87"),
   414 => (x"e6",x"c2",x"87",x"f8"),
   415 => (x"c2",x"4c",x"bf",x"ea"),
   416 => (x"c2",x"5c",x"d3",x"eb"),
   417 => (x"bf",x"97",x"cf",x"df"),
   418 => (x"c2",x"31",x"c8",x"49"),
   419 => (x"bf",x"97",x"ce",x"df"),
   420 => (x"c2",x"49",x"a1",x"4a"),
   421 => (x"bf",x"97",x"d0",x"df"),
   422 => (x"72",x"32",x"d0",x"4a"),
   423 => (x"df",x"c2",x"49",x"a1"),
   424 => (x"4a",x"bf",x"97",x"d1"),
   425 => (x"a1",x"72",x"32",x"d8"),
   426 => (x"91",x"66",x"c4",x"49"),
   427 => (x"bf",x"ff",x"ea",x"c2"),
   428 => (x"c7",x"eb",x"c2",x"81"),
   429 => (x"d7",x"df",x"c2",x"59"),
   430 => (x"c8",x"4a",x"bf",x"97"),
   431 => (x"d6",x"df",x"c2",x"32"),
   432 => (x"a2",x"4b",x"bf",x"97"),
   433 => (x"d8",x"df",x"c2",x"4a"),
   434 => (x"d0",x"4b",x"bf",x"97"),
   435 => (x"4a",x"a2",x"73",x"33"),
   436 => (x"97",x"d9",x"df",x"c2"),
   437 => (x"9b",x"cf",x"4b",x"bf"),
   438 => (x"a2",x"73",x"33",x"d8"),
   439 => (x"cb",x"eb",x"c2",x"4a"),
   440 => (x"c7",x"eb",x"c2",x"5a"),
   441 => (x"8a",x"c2",x"4a",x"bf"),
   442 => (x"eb",x"c2",x"92",x"74"),
   443 => (x"a1",x"72",x"48",x"cb"),
   444 => (x"87",x"ca",x"c1",x"78"),
   445 => (x"97",x"fc",x"de",x"c2"),
   446 => (x"31",x"c8",x"49",x"bf"),
   447 => (x"97",x"fb",x"de",x"c2"),
   448 => (x"49",x"a1",x"4a",x"bf"),
   449 => (x"59",x"fa",x"e6",x"c2"),
   450 => (x"bf",x"f6",x"e6",x"c2"),
   451 => (x"c7",x"31",x"c5",x"49"),
   452 => (x"29",x"c9",x"81",x"ff"),
   453 => (x"59",x"d3",x"eb",x"c2"),
   454 => (x"97",x"c1",x"df",x"c2"),
   455 => (x"32",x"c8",x"4a",x"bf"),
   456 => (x"97",x"c0",x"df",x"c2"),
   457 => (x"4a",x"a2",x"4b",x"bf"),
   458 => (x"6e",x"92",x"66",x"c4"),
   459 => (x"cf",x"eb",x"c2",x"82"),
   460 => (x"c7",x"eb",x"c2",x"5a"),
   461 => (x"c2",x"78",x"c0",x"48"),
   462 => (x"72",x"48",x"c3",x"eb"),
   463 => (x"eb",x"c2",x"78",x"a1"),
   464 => (x"eb",x"c2",x"48",x"d3"),
   465 => (x"c2",x"78",x"bf",x"c7"),
   466 => (x"c2",x"48",x"d7",x"eb"),
   467 => (x"78",x"bf",x"cb",x"eb"),
   468 => (x"bf",x"f2",x"e6",x"c2"),
   469 => (x"87",x"c9",x"c0",x"02"),
   470 => (x"30",x"c4",x"48",x"74"),
   471 => (x"c9",x"c0",x"7e",x"70"),
   472 => (x"cf",x"eb",x"c2",x"87"),
   473 => (x"30",x"c4",x"48",x"bf"),
   474 => (x"e6",x"c2",x"7e",x"70"),
   475 => (x"78",x"6e",x"48",x"f6"),
   476 => (x"8e",x"f8",x"48",x"c1"),
   477 => (x"4c",x"26",x"4d",x"26"),
   478 => (x"4f",x"26",x"4b",x"26"),
   479 => (x"5c",x"5b",x"5e",x"0e"),
   480 => (x"4a",x"71",x"0e",x"5d"),
   481 => (x"bf",x"f2",x"e6",x"c2"),
   482 => (x"72",x"87",x"cb",x"02"),
   483 => (x"72",x"2b",x"c7",x"4b"),
   484 => (x"9c",x"ff",x"c1",x"4c"),
   485 => (x"4b",x"72",x"87",x"c9"),
   486 => (x"4c",x"72",x"2b",x"c8"),
   487 => (x"c2",x"9c",x"ff",x"c3"),
   488 => (x"83",x"bf",x"ff",x"ea"),
   489 => (x"bf",x"c3",x"f2",x"c0"),
   490 => (x"87",x"d9",x"02",x"ab"),
   491 => (x"5b",x"c7",x"f2",x"c0"),
   492 => (x"1e",x"ea",x"de",x"c2"),
   493 => (x"fd",x"f0",x"49",x"73"),
   494 => (x"70",x"86",x"c4",x"87"),
   495 => (x"87",x"c5",x"05",x"98"),
   496 => (x"e6",x"c0",x"48",x"c0"),
   497 => (x"f2",x"e6",x"c2",x"87"),
   498 => (x"87",x"d2",x"02",x"bf"),
   499 => (x"91",x"c4",x"49",x"74"),
   500 => (x"81",x"ea",x"de",x"c2"),
   501 => (x"ff",x"cf",x"4d",x"69"),
   502 => (x"9d",x"ff",x"ff",x"ff"),
   503 => (x"49",x"74",x"87",x"cb"),
   504 => (x"de",x"c2",x"91",x"c2"),
   505 => (x"69",x"9f",x"81",x"ea"),
   506 => (x"fe",x"48",x"75",x"4d"),
   507 => (x"5e",x"0e",x"87",x"c6"),
   508 => (x"0e",x"5d",x"5c",x"5b"),
   509 => (x"c0",x"4d",x"71",x"1e"),
   510 => (x"ca",x"49",x"c1",x"1e"),
   511 => (x"86",x"c4",x"87",x"ee"),
   512 => (x"02",x"9c",x"4c",x"70"),
   513 => (x"c2",x"87",x"c0",x"c1"),
   514 => (x"75",x"4a",x"fa",x"e6"),
   515 => (x"87",x"ff",x"e0",x"49"),
   516 => (x"c0",x"02",x"98",x"70"),
   517 => (x"4a",x"74",x"87",x"f1"),
   518 => (x"4b",x"cb",x"49",x"75"),
   519 => (x"70",x"87",x"e5",x"e1"),
   520 => (x"e2",x"c0",x"02",x"98"),
   521 => (x"74",x"1e",x"c0",x"87"),
   522 => (x"87",x"c7",x"02",x"9c"),
   523 => (x"c0",x"48",x"a6",x"c4"),
   524 => (x"c4",x"87",x"c5",x"78"),
   525 => (x"78",x"c1",x"48",x"a6"),
   526 => (x"c9",x"49",x"66",x"c4"),
   527 => (x"86",x"c4",x"87",x"ee"),
   528 => (x"05",x"9c",x"4c",x"70"),
   529 => (x"74",x"87",x"c0",x"ff"),
   530 => (x"e7",x"fc",x"26",x"48"),
   531 => (x"5b",x"5e",x"0e",x"87"),
   532 => (x"1e",x"0e",x"5d",x"5c"),
   533 => (x"05",x"9b",x"4b",x"71"),
   534 => (x"48",x"c0",x"87",x"c5"),
   535 => (x"c8",x"87",x"e5",x"c1"),
   536 => (x"7d",x"c0",x"4d",x"a3"),
   537 => (x"c7",x"02",x"66",x"d4"),
   538 => (x"97",x"66",x"d4",x"87"),
   539 => (x"87",x"c5",x"05",x"bf"),
   540 => (x"cf",x"c1",x"48",x"c0"),
   541 => (x"49",x"66",x"d4",x"87"),
   542 => (x"70",x"87",x"f3",x"fd"),
   543 => (x"c1",x"02",x"9c",x"4c"),
   544 => (x"a4",x"dc",x"87",x"c0"),
   545 => (x"da",x"7d",x"69",x"49"),
   546 => (x"a3",x"c4",x"49",x"a4"),
   547 => (x"7a",x"69",x"9f",x"4a"),
   548 => (x"bf",x"f2",x"e6",x"c2"),
   549 => (x"d4",x"87",x"d2",x"02"),
   550 => (x"69",x"9f",x"49",x"a4"),
   551 => (x"ff",x"ff",x"c0",x"49"),
   552 => (x"d0",x"48",x"71",x"99"),
   553 => (x"c2",x"7e",x"70",x"30"),
   554 => (x"6e",x"7e",x"c0",x"87"),
   555 => (x"80",x"6a",x"48",x"49"),
   556 => (x"7b",x"c0",x"7a",x"70"),
   557 => (x"6a",x"49",x"a3",x"cc"),
   558 => (x"49",x"a3",x"d0",x"79"),
   559 => (x"48",x"74",x"79",x"c0"),
   560 => (x"48",x"c0",x"87",x"c2"),
   561 => (x"87",x"ec",x"fa",x"26"),
   562 => (x"5c",x"5b",x"5e",x"0e"),
   563 => (x"4c",x"71",x"0e",x"5d"),
   564 => (x"48",x"c3",x"f2",x"c0"),
   565 => (x"9c",x"74",x"78",x"ff"),
   566 => (x"87",x"ca",x"c1",x"02"),
   567 => (x"69",x"49",x"a4",x"c8"),
   568 => (x"87",x"c2",x"c1",x"02"),
   569 => (x"6c",x"4a",x"66",x"d0"),
   570 => (x"a6",x"d4",x"82",x"49"),
   571 => (x"4d",x"66",x"d0",x"5a"),
   572 => (x"ee",x"e6",x"c2",x"b9"),
   573 => (x"ba",x"ff",x"4a",x"bf"),
   574 => (x"99",x"71",x"99",x"72"),
   575 => (x"87",x"e4",x"c0",x"02"),
   576 => (x"6b",x"4b",x"a4",x"c4"),
   577 => (x"87",x"f4",x"f9",x"49"),
   578 => (x"e6",x"c2",x"7b",x"70"),
   579 => (x"6c",x"49",x"bf",x"ea"),
   580 => (x"75",x"7c",x"71",x"81"),
   581 => (x"ee",x"e6",x"c2",x"b9"),
   582 => (x"ba",x"ff",x"4a",x"bf"),
   583 => (x"99",x"71",x"99",x"72"),
   584 => (x"87",x"dc",x"ff",x"05"),
   585 => (x"cb",x"f9",x"7c",x"75"),
   586 => (x"1e",x"73",x"1e",x"87"),
   587 => (x"02",x"9b",x"4b",x"71"),
   588 => (x"a3",x"c8",x"87",x"c7"),
   589 => (x"c5",x"05",x"69",x"49"),
   590 => (x"c0",x"48",x"c0",x"87"),
   591 => (x"eb",x"c2",x"87",x"eb"),
   592 => (x"c4",x"4a",x"bf",x"c3"),
   593 => (x"49",x"69",x"49",x"a3"),
   594 => (x"e6",x"c2",x"89",x"c2"),
   595 => (x"71",x"91",x"bf",x"ea"),
   596 => (x"e6",x"c2",x"4a",x"a2"),
   597 => (x"6b",x"49",x"bf",x"ee"),
   598 => (x"4a",x"a2",x"71",x"99"),
   599 => (x"72",x"1e",x"66",x"c8"),
   600 => (x"87",x"d2",x"ea",x"49"),
   601 => (x"49",x"70",x"86",x"c4"),
   602 => (x"87",x"cc",x"f8",x"48"),
   603 => (x"71",x"1e",x"73",x"1e"),
   604 => (x"c7",x"02",x"9b",x"4b"),
   605 => (x"49",x"a3",x"c8",x"87"),
   606 => (x"87",x"c5",x"05",x"69"),
   607 => (x"eb",x"c0",x"48",x"c0"),
   608 => (x"c3",x"eb",x"c2",x"87"),
   609 => (x"a3",x"c4",x"4a",x"bf"),
   610 => (x"c2",x"49",x"69",x"49"),
   611 => (x"ea",x"e6",x"c2",x"89"),
   612 => (x"a2",x"71",x"91",x"bf"),
   613 => (x"ee",x"e6",x"c2",x"4a"),
   614 => (x"99",x"6b",x"49",x"bf"),
   615 => (x"c8",x"4a",x"a2",x"71"),
   616 => (x"49",x"72",x"1e",x"66"),
   617 => (x"c4",x"87",x"c5",x"e6"),
   618 => (x"48",x"49",x"70",x"86"),
   619 => (x"0e",x"87",x"c9",x"f7"),
   620 => (x"5d",x"5c",x"5b",x"5e"),
   621 => (x"4b",x"71",x"1e",x"0e"),
   622 => (x"c9",x"4c",x"66",x"d4"),
   623 => (x"02",x"9b",x"73",x"2c"),
   624 => (x"c8",x"87",x"cf",x"c1"),
   625 => (x"02",x"69",x"49",x"a3"),
   626 => (x"d0",x"87",x"c7",x"c1"),
   627 => (x"66",x"d4",x"4d",x"a3"),
   628 => (x"ee",x"e6",x"c2",x"7d"),
   629 => (x"b9",x"ff",x"49",x"bf"),
   630 => (x"7e",x"99",x"4a",x"6b"),
   631 => (x"cd",x"03",x"ac",x"71"),
   632 => (x"7d",x"7b",x"c0",x"87"),
   633 => (x"c4",x"4a",x"a3",x"cc"),
   634 => (x"79",x"6a",x"49",x"a3"),
   635 => (x"8c",x"72",x"87",x"c2"),
   636 => (x"dd",x"02",x"9c",x"74"),
   637 => (x"73",x"1e",x"49",x"87"),
   638 => (x"87",x"cc",x"fb",x"49"),
   639 => (x"66",x"d4",x"86",x"c4"),
   640 => (x"99",x"ff",x"c7",x"49"),
   641 => (x"c2",x"87",x"cb",x"02"),
   642 => (x"73",x"1e",x"ea",x"de"),
   643 => (x"87",x"d9",x"fc",x"49"),
   644 => (x"f5",x"26",x"86",x"c4"),
   645 => (x"73",x"1e",x"87",x"de"),
   646 => (x"9b",x"4b",x"71",x"1e"),
   647 => (x"87",x"e4",x"c0",x"02"),
   648 => (x"5b",x"d7",x"eb",x"c2"),
   649 => (x"8a",x"c2",x"4a",x"73"),
   650 => (x"bf",x"ea",x"e6",x"c2"),
   651 => (x"eb",x"c2",x"92",x"49"),
   652 => (x"72",x"48",x"bf",x"c3"),
   653 => (x"db",x"eb",x"c2",x"80"),
   654 => (x"c4",x"48",x"71",x"58"),
   655 => (x"fa",x"e6",x"c2",x"30"),
   656 => (x"87",x"ed",x"c0",x"58"),
   657 => (x"48",x"d3",x"eb",x"c2"),
   658 => (x"bf",x"c7",x"eb",x"c2"),
   659 => (x"d7",x"eb",x"c2",x"78"),
   660 => (x"cb",x"eb",x"c2",x"48"),
   661 => (x"e6",x"c2",x"78",x"bf"),
   662 => (x"c9",x"02",x"bf",x"f2"),
   663 => (x"ea",x"e6",x"c2",x"87"),
   664 => (x"31",x"c4",x"49",x"bf"),
   665 => (x"eb",x"c2",x"87",x"c7"),
   666 => (x"c4",x"49",x"bf",x"cf"),
   667 => (x"fa",x"e6",x"c2",x"31"),
   668 => (x"87",x"c4",x"f4",x"59"),
   669 => (x"5c",x"5b",x"5e",x"0e"),
   670 => (x"c0",x"4a",x"71",x"0e"),
   671 => (x"02",x"9a",x"72",x"4b"),
   672 => (x"da",x"87",x"e1",x"c0"),
   673 => (x"69",x"9f",x"49",x"a2"),
   674 => (x"f2",x"e6",x"c2",x"4b"),
   675 => (x"87",x"cf",x"02",x"bf"),
   676 => (x"9f",x"49",x"a2",x"d4"),
   677 => (x"c0",x"4c",x"49",x"69"),
   678 => (x"d0",x"9c",x"ff",x"ff"),
   679 => (x"c0",x"87",x"c2",x"34"),
   680 => (x"b3",x"49",x"74",x"4c"),
   681 => (x"ed",x"fd",x"49",x"73"),
   682 => (x"87",x"ca",x"f3",x"87"),
   683 => (x"5c",x"5b",x"5e",x"0e"),
   684 => (x"86",x"f4",x"0e",x"5d"),
   685 => (x"7e",x"c0",x"4a",x"71"),
   686 => (x"d8",x"02",x"9a",x"72"),
   687 => (x"e6",x"de",x"c2",x"87"),
   688 => (x"c2",x"78",x"c0",x"48"),
   689 => (x"c2",x"48",x"de",x"de"),
   690 => (x"78",x"bf",x"d7",x"eb"),
   691 => (x"48",x"e2",x"de",x"c2"),
   692 => (x"bf",x"d3",x"eb",x"c2"),
   693 => (x"c7",x"e7",x"c2",x"78"),
   694 => (x"c2",x"50",x"c0",x"48"),
   695 => (x"49",x"bf",x"f6",x"e6"),
   696 => (x"bf",x"e6",x"de",x"c2"),
   697 => (x"03",x"aa",x"71",x"4a"),
   698 => (x"72",x"87",x"ff",x"c3"),
   699 => (x"05",x"99",x"cf",x"49"),
   700 => (x"c2",x"87",x"e0",x"c0"),
   701 => (x"c2",x"1e",x"ea",x"de"),
   702 => (x"49",x"bf",x"de",x"de"),
   703 => (x"48",x"de",x"de",x"c2"),
   704 => (x"71",x"78",x"a1",x"c1"),
   705 => (x"c4",x"87",x"ef",x"e3"),
   706 => (x"ff",x"f1",x"c0",x"86"),
   707 => (x"ea",x"de",x"c2",x"48"),
   708 => (x"c0",x"87",x"cc",x"78"),
   709 => (x"48",x"bf",x"ff",x"f1"),
   710 => (x"c0",x"80",x"e0",x"c0"),
   711 => (x"c2",x"58",x"c3",x"f2"),
   712 => (x"48",x"bf",x"e6",x"de"),
   713 => (x"de",x"c2",x"80",x"c1"),
   714 => (x"7f",x"27",x"58",x"ea"),
   715 => (x"bf",x"00",x"00",x"0c"),
   716 => (x"9d",x"4d",x"bf",x"97"),
   717 => (x"87",x"e2",x"c2",x"02"),
   718 => (x"02",x"ad",x"e5",x"c3"),
   719 => (x"c0",x"87",x"db",x"c2"),
   720 => (x"4b",x"bf",x"ff",x"f1"),
   721 => (x"11",x"49",x"a3",x"cb"),
   722 => (x"05",x"ac",x"cf",x"4c"),
   723 => (x"75",x"87",x"d2",x"c1"),
   724 => (x"c1",x"99",x"df",x"49"),
   725 => (x"c2",x"91",x"cd",x"89"),
   726 => (x"c1",x"81",x"fa",x"e6"),
   727 => (x"51",x"12",x"4a",x"a3"),
   728 => (x"12",x"4a",x"a3",x"c3"),
   729 => (x"4a",x"a3",x"c5",x"51"),
   730 => (x"a3",x"c7",x"51",x"12"),
   731 => (x"c9",x"51",x"12",x"4a"),
   732 => (x"51",x"12",x"4a",x"a3"),
   733 => (x"12",x"4a",x"a3",x"ce"),
   734 => (x"4a",x"a3",x"d0",x"51"),
   735 => (x"a3",x"d2",x"51",x"12"),
   736 => (x"d4",x"51",x"12",x"4a"),
   737 => (x"51",x"12",x"4a",x"a3"),
   738 => (x"12",x"4a",x"a3",x"d6"),
   739 => (x"4a",x"a3",x"d8",x"51"),
   740 => (x"a3",x"dc",x"51",x"12"),
   741 => (x"de",x"51",x"12",x"4a"),
   742 => (x"51",x"12",x"4a",x"a3"),
   743 => (x"f9",x"c0",x"7e",x"c1"),
   744 => (x"c8",x"49",x"74",x"87"),
   745 => (x"ea",x"c0",x"05",x"99"),
   746 => (x"d0",x"49",x"74",x"87"),
   747 => (x"87",x"d0",x"05",x"99"),
   748 => (x"c0",x"02",x"66",x"dc"),
   749 => (x"49",x"73",x"87",x"ca"),
   750 => (x"70",x"0f",x"66",x"dc"),
   751 => (x"87",x"d3",x"02",x"98"),
   752 => (x"c6",x"c0",x"05",x"6e"),
   753 => (x"fa",x"e6",x"c2",x"87"),
   754 => (x"c0",x"50",x"c0",x"48"),
   755 => (x"48",x"bf",x"ff",x"f1"),
   756 => (x"c2",x"87",x"e7",x"c2"),
   757 => (x"c0",x"48",x"c7",x"e7"),
   758 => (x"e6",x"c2",x"7e",x"50"),
   759 => (x"c2",x"49",x"bf",x"f6"),
   760 => (x"4a",x"bf",x"e6",x"de"),
   761 => (x"fc",x"04",x"aa",x"71"),
   762 => (x"eb",x"c2",x"87",x"c1"),
   763 => (x"c0",x"05",x"bf",x"d7"),
   764 => (x"e6",x"c2",x"87",x"c8"),
   765 => (x"c1",x"02",x"bf",x"f2"),
   766 => (x"f2",x"c0",x"87",x"fe"),
   767 => (x"78",x"ff",x"48",x"c3"),
   768 => (x"bf",x"e2",x"de",x"c2"),
   769 => (x"87",x"f4",x"ed",x"49"),
   770 => (x"de",x"c2",x"49",x"70"),
   771 => (x"a6",x"c4",x"59",x"e6"),
   772 => (x"e2",x"de",x"c2",x"48"),
   773 => (x"e6",x"c2",x"78",x"bf"),
   774 => (x"c0",x"02",x"bf",x"f2"),
   775 => (x"66",x"c4",x"87",x"d8"),
   776 => (x"ff",x"ff",x"cf",x"49"),
   777 => (x"a9",x"99",x"f8",x"ff"),
   778 => (x"87",x"c5",x"c0",x"02"),
   779 => (x"e1",x"c0",x"4d",x"c0"),
   780 => (x"c0",x"4d",x"c1",x"87"),
   781 => (x"66",x"c4",x"87",x"dc"),
   782 => (x"f8",x"ff",x"cf",x"49"),
   783 => (x"c0",x"02",x"a9",x"99"),
   784 => (x"a6",x"c8",x"87",x"c8"),
   785 => (x"c0",x"78",x"c0",x"48"),
   786 => (x"a6",x"c8",x"87",x"c5"),
   787 => (x"c8",x"78",x"c1",x"48"),
   788 => (x"9d",x"75",x"4d",x"66"),
   789 => (x"87",x"e0",x"c0",x"05"),
   790 => (x"c2",x"49",x"66",x"c4"),
   791 => (x"ea",x"e6",x"c2",x"89"),
   792 => (x"c2",x"91",x"4a",x"bf"),
   793 => (x"4a",x"bf",x"c3",x"eb"),
   794 => (x"48",x"de",x"de",x"c2"),
   795 => (x"c2",x"78",x"a1",x"72"),
   796 => (x"c0",x"48",x"e6",x"de"),
   797 => (x"87",x"e3",x"f9",x"78"),
   798 => (x"8e",x"f4",x"48",x"c0"),
   799 => (x"00",x"87",x"f5",x"eb"),
   800 => (x"ff",x"00",x"00",x"00"),
   801 => (x"8f",x"ff",x"ff",x"ff"),
   802 => (x"98",x"00",x"00",x"0c"),
   803 => (x"46",x"00",x"00",x"0c"),
   804 => (x"32",x"33",x"54",x"41"),
   805 => (x"00",x"20",x"20",x"20"),
   806 => (x"31",x"54",x"41",x"46"),
   807 => (x"20",x"20",x"20",x"36"),
   808 => (x"d4",x"ff",x"1e",x"00"),
   809 => (x"78",x"ff",x"c3",x"48"),
   810 => (x"4f",x"26",x"48",x"68"),
   811 => (x"48",x"d4",x"ff",x"1e"),
   812 => (x"ff",x"78",x"ff",x"c3"),
   813 => (x"e1",x"c8",x"48",x"d0"),
   814 => (x"48",x"d4",x"ff",x"78"),
   815 => (x"eb",x"c2",x"78",x"d4"),
   816 => (x"d4",x"ff",x"48",x"db"),
   817 => (x"4f",x"26",x"50",x"bf"),
   818 => (x"48",x"d0",x"ff",x"1e"),
   819 => (x"26",x"78",x"e0",x"c0"),
   820 => (x"cc",x"ff",x"1e",x"4f"),
   821 => (x"99",x"49",x"70",x"87"),
   822 => (x"c0",x"87",x"c6",x"02"),
   823 => (x"f1",x"05",x"a9",x"fb"),
   824 => (x"26",x"48",x"71",x"87"),
   825 => (x"5b",x"5e",x"0e",x"4f"),
   826 => (x"4b",x"71",x"0e",x"5c"),
   827 => (x"f0",x"fe",x"4c",x"c0"),
   828 => (x"99",x"49",x"70",x"87"),
   829 => (x"87",x"f9",x"c0",x"02"),
   830 => (x"02",x"a9",x"ec",x"c0"),
   831 => (x"c0",x"87",x"f2",x"c0"),
   832 => (x"c0",x"02",x"a9",x"fb"),
   833 => (x"66",x"cc",x"87",x"eb"),
   834 => (x"c7",x"03",x"ac",x"b7"),
   835 => (x"02",x"66",x"d0",x"87"),
   836 => (x"53",x"71",x"87",x"c2"),
   837 => (x"c2",x"02",x"99",x"71"),
   838 => (x"fe",x"84",x"c1",x"87"),
   839 => (x"49",x"70",x"87",x"c3"),
   840 => (x"87",x"cd",x"02",x"99"),
   841 => (x"02",x"a9",x"ec",x"c0"),
   842 => (x"fb",x"c0",x"87",x"c7"),
   843 => (x"d5",x"ff",x"05",x"a9"),
   844 => (x"02",x"66",x"d0",x"87"),
   845 => (x"97",x"c0",x"87",x"c3"),
   846 => (x"a9",x"ec",x"c0",x"7b"),
   847 => (x"74",x"87",x"c4",x"05"),
   848 => (x"74",x"87",x"c5",x"4a"),
   849 => (x"8a",x"0a",x"c0",x"4a"),
   850 => (x"87",x"c2",x"48",x"72"),
   851 => (x"4c",x"26",x"4d",x"26"),
   852 => (x"4f",x"26",x"4b",x"26"),
   853 => (x"87",x"c9",x"fd",x"1e"),
   854 => (x"f0",x"c0",x"49",x"70"),
   855 => (x"ca",x"04",x"a9",x"b7"),
   856 => (x"b7",x"f9",x"c0",x"87"),
   857 => (x"87",x"c3",x"01",x"a9"),
   858 => (x"c1",x"89",x"f0",x"c0"),
   859 => (x"04",x"a9",x"b7",x"c1"),
   860 => (x"da",x"c1",x"87",x"ca"),
   861 => (x"c3",x"01",x"a9",x"b7"),
   862 => (x"89",x"f7",x"c0",x"87"),
   863 => (x"4f",x"26",x"48",x"71"),
   864 => (x"5c",x"5b",x"5e",x"0e"),
   865 => (x"ff",x"4a",x"71",x"0e"),
   866 => (x"49",x"72",x"4c",x"d4"),
   867 => (x"70",x"87",x"ea",x"c0"),
   868 => (x"c2",x"02",x"9b",x"4b"),
   869 => (x"ff",x"8b",x"c1",x"87"),
   870 => (x"c5",x"c8",x"48",x"d0"),
   871 => (x"7c",x"d5",x"c1",x"78"),
   872 => (x"31",x"c6",x"49",x"73"),
   873 => (x"97",x"db",x"dc",x"c2"),
   874 => (x"71",x"48",x"4a",x"bf"),
   875 => (x"ff",x"7c",x"70",x"b0"),
   876 => (x"78",x"c4",x"48",x"d0"),
   877 => (x"d5",x"fe",x"48",x"73"),
   878 => (x"5b",x"5e",x"0e",x"87"),
   879 => (x"f8",x"0e",x"5d",x"5c"),
   880 => (x"c0",x"4c",x"71",x"86"),
   881 => (x"87",x"e4",x"fb",x"7e"),
   882 => (x"f9",x"c0",x"4b",x"c0"),
   883 => (x"49",x"bf",x"97",x"e6"),
   884 => (x"cf",x"04",x"a9",x"c0"),
   885 => (x"87",x"f9",x"fb",x"87"),
   886 => (x"f9",x"c0",x"83",x"c1"),
   887 => (x"49",x"bf",x"97",x"e6"),
   888 => (x"87",x"f1",x"06",x"ab"),
   889 => (x"97",x"e6",x"f9",x"c0"),
   890 => (x"87",x"cf",x"02",x"bf"),
   891 => (x"70",x"87",x"f2",x"fa"),
   892 => (x"c6",x"02",x"99",x"49"),
   893 => (x"a9",x"ec",x"c0",x"87"),
   894 => (x"c0",x"87",x"f1",x"05"),
   895 => (x"87",x"e1",x"fa",x"4b"),
   896 => (x"dc",x"fa",x"4d",x"70"),
   897 => (x"58",x"a6",x"c8",x"87"),
   898 => (x"70",x"87",x"d6",x"fa"),
   899 => (x"c8",x"83",x"c1",x"4a"),
   900 => (x"69",x"97",x"49",x"a4"),
   901 => (x"c7",x"02",x"ad",x"49"),
   902 => (x"ad",x"ff",x"c0",x"87"),
   903 => (x"87",x"e7",x"c0",x"05"),
   904 => (x"97",x"49",x"a4",x"c9"),
   905 => (x"66",x"c4",x"49",x"69"),
   906 => (x"87",x"c7",x"02",x"a9"),
   907 => (x"a8",x"ff",x"c0",x"48"),
   908 => (x"ca",x"87",x"d4",x"05"),
   909 => (x"69",x"97",x"49",x"a4"),
   910 => (x"c6",x"02",x"aa",x"49"),
   911 => (x"aa",x"ff",x"c0",x"87"),
   912 => (x"c1",x"87",x"c4",x"05"),
   913 => (x"c0",x"87",x"d0",x"7e"),
   914 => (x"c6",x"02",x"ad",x"ec"),
   915 => (x"ad",x"fb",x"c0",x"87"),
   916 => (x"c0",x"87",x"c4",x"05"),
   917 => (x"6e",x"7e",x"c1",x"4b"),
   918 => (x"87",x"e1",x"fe",x"02"),
   919 => (x"73",x"87",x"e9",x"f9"),
   920 => (x"fb",x"8e",x"f8",x"48"),
   921 => (x"0e",x"00",x"87",x"e6"),
   922 => (x"5d",x"5c",x"5b",x"5e"),
   923 => (x"4b",x"71",x"1e",x"0e"),
   924 => (x"ab",x"4d",x"4c",x"c0"),
   925 => (x"87",x"e8",x"c0",x"04"),
   926 => (x"1e",x"f9",x"f6",x"c0"),
   927 => (x"c4",x"02",x"9d",x"75"),
   928 => (x"c2",x"4a",x"c0",x"87"),
   929 => (x"72",x"4a",x"c1",x"87"),
   930 => (x"87",x"e0",x"f0",x"49"),
   931 => (x"7e",x"70",x"86",x"c4"),
   932 => (x"05",x"6e",x"84",x"c1"),
   933 => (x"4c",x"73",x"87",x"c2"),
   934 => (x"ac",x"73",x"85",x"c1"),
   935 => (x"87",x"d8",x"ff",x"06"),
   936 => (x"26",x"26",x"48",x"6e"),
   937 => (x"26",x"4c",x"26",x"4d"),
   938 => (x"0e",x"4f",x"26",x"4b"),
   939 => (x"5d",x"5c",x"5b",x"5e"),
   940 => (x"4c",x"71",x"1e",x"0e"),
   941 => (x"c2",x"91",x"de",x"49"),
   942 => (x"71",x"4d",x"f5",x"eb"),
   943 => (x"02",x"6d",x"97",x"85"),
   944 => (x"c2",x"87",x"dd",x"c1"),
   945 => (x"4a",x"bf",x"e0",x"eb"),
   946 => (x"49",x"72",x"82",x"74"),
   947 => (x"70",x"87",x"d8",x"fe"),
   948 => (x"c0",x"02",x"6e",x"7e"),
   949 => (x"eb",x"c2",x"87",x"f3"),
   950 => (x"4a",x"6e",x"4b",x"e8"),
   951 => (x"c7",x"ff",x"49",x"cb"),
   952 => (x"4b",x"74",x"87",x"c6"),
   953 => (x"dd",x"c1",x"93",x"cb"),
   954 => (x"83",x"c4",x"83",x"e7"),
   955 => (x"7b",x"e4",x"fc",x"c0"),
   956 => (x"c4",x"c1",x"49",x"74"),
   957 => (x"7b",x"75",x"87",x"dc"),
   958 => (x"97",x"f4",x"eb",x"c2"),
   959 => (x"c2",x"1e",x"49",x"bf"),
   960 => (x"c1",x"49",x"e8",x"eb"),
   961 => (x"c4",x"87",x"d6",x"df"),
   962 => (x"c1",x"49",x"74",x"86"),
   963 => (x"c0",x"87",x"c3",x"c4"),
   964 => (x"e2",x"c5",x"c1",x"49"),
   965 => (x"dc",x"eb",x"c2",x"87"),
   966 => (x"c1",x"78",x"c0",x"48"),
   967 => (x"87",x"f9",x"dc",x"49"),
   968 => (x"87",x"ff",x"fd",x"26"),
   969 => (x"64",x"61",x"6f",x"4c"),
   970 => (x"2e",x"67",x"6e",x"69"),
   971 => (x"0e",x"00",x"2e",x"2e"),
   972 => (x"0e",x"5c",x"5b",x"5e"),
   973 => (x"c2",x"4a",x"4b",x"71"),
   974 => (x"82",x"bf",x"e0",x"eb"),
   975 => (x"e6",x"fc",x"49",x"72"),
   976 => (x"9c",x"4c",x"70",x"87"),
   977 => (x"49",x"87",x"c4",x"02"),
   978 => (x"c2",x"87",x"e9",x"ec"),
   979 => (x"c0",x"48",x"e0",x"eb"),
   980 => (x"dc",x"49",x"c1",x"78"),
   981 => (x"cc",x"fd",x"87",x"c3"),
   982 => (x"5b",x"5e",x"0e",x"87"),
   983 => (x"f4",x"0e",x"5d",x"5c"),
   984 => (x"ea",x"de",x"c2",x"86"),
   985 => (x"c4",x"4c",x"c0",x"4d"),
   986 => (x"78",x"c0",x"48",x"a6"),
   987 => (x"bf",x"e0",x"eb",x"c2"),
   988 => (x"06",x"a9",x"c0",x"49"),
   989 => (x"c2",x"87",x"c1",x"c1"),
   990 => (x"98",x"48",x"ea",x"de"),
   991 => (x"87",x"f8",x"c0",x"02"),
   992 => (x"1e",x"f9",x"f6",x"c0"),
   993 => (x"c7",x"02",x"66",x"c8"),
   994 => (x"48",x"a6",x"c4",x"87"),
   995 => (x"87",x"c5",x"78",x"c0"),
   996 => (x"c1",x"48",x"a6",x"c4"),
   997 => (x"49",x"66",x"c4",x"78"),
   998 => (x"c4",x"87",x"d1",x"ec"),
   999 => (x"c1",x"4d",x"70",x"86"),
  1000 => (x"48",x"66",x"c4",x"84"),
  1001 => (x"a6",x"c8",x"80",x"c1"),
  1002 => (x"e0",x"eb",x"c2",x"58"),
  1003 => (x"03",x"ac",x"49",x"bf"),
  1004 => (x"9d",x"75",x"87",x"c6"),
  1005 => (x"87",x"c8",x"ff",x"05"),
  1006 => (x"9d",x"75",x"4c",x"c0"),
  1007 => (x"87",x"e0",x"c3",x"02"),
  1008 => (x"1e",x"f9",x"f6",x"c0"),
  1009 => (x"c7",x"02",x"66",x"c8"),
  1010 => (x"48",x"a6",x"cc",x"87"),
  1011 => (x"87",x"c5",x"78",x"c0"),
  1012 => (x"c1",x"48",x"a6",x"cc"),
  1013 => (x"49",x"66",x"cc",x"78"),
  1014 => (x"c4",x"87",x"d1",x"eb"),
  1015 => (x"6e",x"7e",x"70",x"86"),
  1016 => (x"87",x"e9",x"c2",x"02"),
  1017 => (x"81",x"cb",x"49",x"6e"),
  1018 => (x"d0",x"49",x"69",x"97"),
  1019 => (x"d6",x"c1",x"02",x"99"),
  1020 => (x"ef",x"fc",x"c0",x"87"),
  1021 => (x"cb",x"49",x"74",x"4a"),
  1022 => (x"e7",x"dd",x"c1",x"91"),
  1023 => (x"c8",x"79",x"72",x"81"),
  1024 => (x"51",x"ff",x"c3",x"81"),
  1025 => (x"91",x"de",x"49",x"74"),
  1026 => (x"4d",x"f5",x"eb",x"c2"),
  1027 => (x"c1",x"c2",x"85",x"71"),
  1028 => (x"a5",x"c1",x"7d",x"97"),
  1029 => (x"51",x"e0",x"c0",x"49"),
  1030 => (x"97",x"fa",x"e6",x"c2"),
  1031 => (x"87",x"d2",x"02",x"bf"),
  1032 => (x"a5",x"c2",x"84",x"c1"),
  1033 => (x"fa",x"e6",x"c2",x"4b"),
  1034 => (x"ff",x"49",x"db",x"4a"),
  1035 => (x"c1",x"87",x"f9",x"c1"),
  1036 => (x"a5",x"cd",x"87",x"db"),
  1037 => (x"c1",x"51",x"c0",x"49"),
  1038 => (x"4b",x"a5",x"c2",x"84"),
  1039 => (x"49",x"cb",x"4a",x"6e"),
  1040 => (x"87",x"e4",x"c1",x"ff"),
  1041 => (x"c0",x"87",x"c6",x"c1"),
  1042 => (x"74",x"4a",x"eb",x"fa"),
  1043 => (x"c1",x"91",x"cb",x"49"),
  1044 => (x"72",x"81",x"e7",x"dd"),
  1045 => (x"fa",x"e6",x"c2",x"79"),
  1046 => (x"d8",x"02",x"bf",x"97"),
  1047 => (x"de",x"49",x"74",x"87"),
  1048 => (x"c2",x"84",x"c1",x"91"),
  1049 => (x"71",x"4b",x"f5",x"eb"),
  1050 => (x"fa",x"e6",x"c2",x"83"),
  1051 => (x"ff",x"49",x"dd",x"4a"),
  1052 => (x"d8",x"87",x"f5",x"c0"),
  1053 => (x"de",x"4b",x"74",x"87"),
  1054 => (x"f5",x"eb",x"c2",x"93"),
  1055 => (x"49",x"a3",x"cb",x"83"),
  1056 => (x"84",x"c1",x"51",x"c0"),
  1057 => (x"cb",x"4a",x"6e",x"73"),
  1058 => (x"db",x"c0",x"ff",x"49"),
  1059 => (x"48",x"66",x"c4",x"87"),
  1060 => (x"a6",x"c8",x"80",x"c1"),
  1061 => (x"03",x"ac",x"c7",x"58"),
  1062 => (x"6e",x"87",x"c5",x"c0"),
  1063 => (x"87",x"e0",x"fc",x"05"),
  1064 => (x"8e",x"f4",x"48",x"74"),
  1065 => (x"1e",x"87",x"fc",x"f7"),
  1066 => (x"4b",x"71",x"1e",x"73"),
  1067 => (x"c1",x"91",x"cb",x"49"),
  1068 => (x"c8",x"81",x"e7",x"dd"),
  1069 => (x"dc",x"c2",x"4a",x"a1"),
  1070 => (x"50",x"12",x"48",x"db"),
  1071 => (x"c0",x"4a",x"a1",x"c9"),
  1072 => (x"12",x"48",x"e6",x"f9"),
  1073 => (x"c2",x"81",x"ca",x"50"),
  1074 => (x"11",x"48",x"f4",x"eb"),
  1075 => (x"f4",x"eb",x"c2",x"50"),
  1076 => (x"1e",x"49",x"bf",x"97"),
  1077 => (x"d8",x"c1",x"49",x"c0"),
  1078 => (x"eb",x"c2",x"87",x"c3"),
  1079 => (x"78",x"de",x"48",x"dc"),
  1080 => (x"f4",x"d5",x"49",x"c1"),
  1081 => (x"fe",x"f6",x"26",x"87"),
  1082 => (x"4a",x"71",x"1e",x"87"),
  1083 => (x"c1",x"91",x"cb",x"49"),
  1084 => (x"c8",x"81",x"e7",x"dd"),
  1085 => (x"c2",x"48",x"11",x"81"),
  1086 => (x"c2",x"58",x"e0",x"eb"),
  1087 => (x"c0",x"48",x"e0",x"eb"),
  1088 => (x"d5",x"49",x"c1",x"78"),
  1089 => (x"4f",x"26",x"87",x"d3"),
  1090 => (x"c0",x"49",x"c0",x"1e"),
  1091 => (x"26",x"87",x"e8",x"fd"),
  1092 => (x"99",x"71",x"1e",x"4f"),
  1093 => (x"c1",x"87",x"d2",x"02"),
  1094 => (x"c0",x"48",x"fc",x"de"),
  1095 => (x"c1",x"80",x"f7",x"50"),
  1096 => (x"c1",x"40",x"e9",x"c3"),
  1097 => (x"ce",x"78",x"e0",x"dd"),
  1098 => (x"f8",x"de",x"c1",x"87"),
  1099 => (x"d9",x"dd",x"c1",x"48"),
  1100 => (x"c1",x"80",x"fc",x"78"),
  1101 => (x"26",x"78",x"c8",x"c4"),
  1102 => (x"5b",x"5e",x"0e",x"4f"),
  1103 => (x"4c",x"71",x"0e",x"5c"),
  1104 => (x"c1",x"92",x"cb",x"4a"),
  1105 => (x"c8",x"82",x"e7",x"dd"),
  1106 => (x"a2",x"c9",x"49",x"a2"),
  1107 => (x"4b",x"6b",x"97",x"4b"),
  1108 => (x"49",x"69",x"97",x"1e"),
  1109 => (x"12",x"82",x"ca",x"1e"),
  1110 => (x"e3",x"e8",x"c0",x"49"),
  1111 => (x"d3",x"49",x"c0",x"87"),
  1112 => (x"49",x"74",x"87",x"f7"),
  1113 => (x"87",x"ea",x"fa",x"c0"),
  1114 => (x"f8",x"f4",x"8e",x"f8"),
  1115 => (x"1e",x"73",x"1e",x"87"),
  1116 => (x"ff",x"49",x"4b",x"71"),
  1117 => (x"49",x"73",x"87",x"c3"),
  1118 => (x"f4",x"87",x"fe",x"fe"),
  1119 => (x"73",x"1e",x"87",x"e9"),
  1120 => (x"c6",x"4b",x"71",x"1e"),
  1121 => (x"db",x"02",x"4a",x"a3"),
  1122 => (x"02",x"8a",x"c1",x"87"),
  1123 => (x"02",x"8a",x"87",x"d6"),
  1124 => (x"8a",x"87",x"da",x"c1"),
  1125 => (x"87",x"fc",x"c0",x"02"),
  1126 => (x"e1",x"c0",x"02",x"8a"),
  1127 => (x"cb",x"02",x"8a",x"87"),
  1128 => (x"87",x"db",x"c1",x"87"),
  1129 => (x"c0",x"fd",x"49",x"c7"),
  1130 => (x"87",x"de",x"c1",x"87"),
  1131 => (x"bf",x"e0",x"eb",x"c2"),
  1132 => (x"87",x"cb",x"c1",x"02"),
  1133 => (x"c2",x"88",x"c1",x"48"),
  1134 => (x"c1",x"58",x"e4",x"eb"),
  1135 => (x"eb",x"c2",x"87",x"c1"),
  1136 => (x"c0",x"02",x"bf",x"e4"),
  1137 => (x"eb",x"c2",x"87",x"f9"),
  1138 => (x"c1",x"48",x"bf",x"e0"),
  1139 => (x"e4",x"eb",x"c2",x"80"),
  1140 => (x"87",x"eb",x"c0",x"58"),
  1141 => (x"bf",x"e0",x"eb",x"c2"),
  1142 => (x"c2",x"89",x"c6",x"49"),
  1143 => (x"c0",x"59",x"e4",x"eb"),
  1144 => (x"da",x"03",x"a9",x"b7"),
  1145 => (x"e0",x"eb",x"c2",x"87"),
  1146 => (x"d2",x"78",x"c0",x"48"),
  1147 => (x"e4",x"eb",x"c2",x"87"),
  1148 => (x"87",x"cb",x"02",x"bf"),
  1149 => (x"bf",x"e0",x"eb",x"c2"),
  1150 => (x"c2",x"80",x"c6",x"48"),
  1151 => (x"c0",x"58",x"e4",x"eb"),
  1152 => (x"87",x"d5",x"d1",x"49"),
  1153 => (x"f8",x"c0",x"49",x"73"),
  1154 => (x"da",x"f2",x"87",x"c8"),
  1155 => (x"5b",x"5e",x"0e",x"87"),
  1156 => (x"4c",x"71",x"0e",x"5c"),
  1157 => (x"74",x"1e",x"66",x"cc"),
  1158 => (x"c1",x"93",x"cb",x"4b"),
  1159 => (x"c4",x"83",x"e7",x"dd"),
  1160 => (x"49",x"6a",x"4a",x"a3"),
  1161 => (x"87",x"d0",x"fa",x"fe"),
  1162 => (x"7b",x"e7",x"c2",x"c1"),
  1163 => (x"d4",x"49",x"a3",x"c8"),
  1164 => (x"a3",x"c9",x"51",x"66"),
  1165 => (x"51",x"66",x"d8",x"49"),
  1166 => (x"dc",x"49",x"a3",x"ca"),
  1167 => (x"f1",x"26",x"51",x"66"),
  1168 => (x"5e",x"0e",x"87",x"e3"),
  1169 => (x"0e",x"5d",x"5c",x"5b"),
  1170 => (x"d8",x"86",x"d0",x"ff"),
  1171 => (x"a6",x"c4",x"59",x"a6"),
  1172 => (x"c4",x"78",x"c0",x"48"),
  1173 => (x"66",x"c4",x"c1",x"80"),
  1174 => (x"c1",x"80",x"c4",x"78"),
  1175 => (x"c1",x"80",x"c4",x"78"),
  1176 => (x"e4",x"eb",x"c2",x"78"),
  1177 => (x"c2",x"78",x"c1",x"48"),
  1178 => (x"48",x"bf",x"dc",x"eb"),
  1179 => (x"cb",x"05",x"a8",x"de"),
  1180 => (x"87",x"e5",x"f3",x"87"),
  1181 => (x"a6",x"c8",x"49",x"70"),
  1182 => (x"87",x"e6",x"ce",x"59"),
  1183 => (x"e9",x"87",x"ed",x"e8"),
  1184 => (x"dc",x"e8",x"87",x"cf"),
  1185 => (x"c0",x"4c",x"70",x"87"),
  1186 => (x"c1",x"02",x"ac",x"fb"),
  1187 => (x"66",x"d4",x"87",x"d0"),
  1188 => (x"87",x"c2",x"c1",x"05"),
  1189 => (x"c1",x"1e",x"1e",x"c0"),
  1190 => (x"da",x"df",x"c1",x"1e"),
  1191 => (x"fd",x"49",x"c0",x"1e"),
  1192 => (x"d0",x"c1",x"87",x"eb"),
  1193 => (x"82",x"c4",x"4a",x"66"),
  1194 => (x"81",x"c7",x"49",x"6a"),
  1195 => (x"1e",x"c1",x"51",x"74"),
  1196 => (x"49",x"6a",x"1e",x"d8"),
  1197 => (x"ec",x"e8",x"81",x"c8"),
  1198 => (x"c1",x"86",x"d8",x"87"),
  1199 => (x"c0",x"48",x"66",x"c4"),
  1200 => (x"87",x"c7",x"01",x"a8"),
  1201 => (x"c1",x"48",x"a6",x"c4"),
  1202 => (x"c1",x"87",x"ce",x"78"),
  1203 => (x"c1",x"48",x"66",x"c4"),
  1204 => (x"58",x"a6",x"cc",x"88"),
  1205 => (x"f8",x"e7",x"87",x"c3"),
  1206 => (x"48",x"a6",x"cc",x"87"),
  1207 => (x"9c",x"74",x"78",x"c2"),
  1208 => (x"87",x"fa",x"cc",x"02"),
  1209 => (x"c1",x"48",x"66",x"c4"),
  1210 => (x"03",x"a8",x"66",x"c8"),
  1211 => (x"d8",x"87",x"ef",x"cc"),
  1212 => (x"78",x"c0",x"48",x"a6"),
  1213 => (x"78",x"c0",x"80",x"c4"),
  1214 => (x"70",x"87",x"e6",x"e6"),
  1215 => (x"ac",x"d0",x"c1",x"4c"),
  1216 => (x"87",x"d7",x"c2",x"05"),
  1217 => (x"e9",x"7e",x"66",x"dc"),
  1218 => (x"49",x"70",x"87",x"ca"),
  1219 => (x"59",x"a6",x"e0",x"c0"),
  1220 => (x"70",x"87",x"ce",x"e6"),
  1221 => (x"ac",x"ec",x"c0",x"4c"),
  1222 => (x"87",x"ea",x"c1",x"05"),
  1223 => (x"cb",x"49",x"66",x"c4"),
  1224 => (x"66",x"c0",x"c1",x"91"),
  1225 => (x"4a",x"a1",x"c4",x"81"),
  1226 => (x"a1",x"c8",x"4d",x"6a"),
  1227 => (x"52",x"66",x"dc",x"4a"),
  1228 => (x"79",x"e9",x"c3",x"c1"),
  1229 => (x"70",x"87",x"ea",x"e5"),
  1230 => (x"d8",x"02",x"9c",x"4c"),
  1231 => (x"ac",x"fb",x"c0",x"87"),
  1232 => (x"74",x"87",x"d2",x"02"),
  1233 => (x"87",x"d9",x"e5",x"55"),
  1234 => (x"02",x"9c",x"4c",x"70"),
  1235 => (x"fb",x"c0",x"87",x"c7"),
  1236 => (x"ee",x"ff",x"05",x"ac"),
  1237 => (x"55",x"e0",x"c0",x"87"),
  1238 => (x"c0",x"55",x"c1",x"c2"),
  1239 => (x"66",x"d4",x"7d",x"97"),
  1240 => (x"05",x"a9",x"6e",x"49"),
  1241 => (x"66",x"c4",x"87",x"db"),
  1242 => (x"a8",x"66",x"c8",x"48"),
  1243 => (x"c4",x"87",x"ca",x"04"),
  1244 => (x"80",x"c1",x"48",x"66"),
  1245 => (x"c8",x"58",x"a6",x"c8"),
  1246 => (x"48",x"66",x"c8",x"87"),
  1247 => (x"a6",x"cc",x"88",x"c1"),
  1248 => (x"87",x"dd",x"e4",x"58"),
  1249 => (x"d0",x"c1",x"4c",x"70"),
  1250 => (x"87",x"c8",x"05",x"ac"),
  1251 => (x"c1",x"48",x"66",x"d0"),
  1252 => (x"58",x"a6",x"d4",x"80"),
  1253 => (x"02",x"ac",x"d0",x"c1"),
  1254 => (x"c0",x"87",x"e9",x"fd"),
  1255 => (x"d4",x"48",x"a6",x"e0"),
  1256 => (x"66",x"dc",x"78",x"66"),
  1257 => (x"66",x"e0",x"c0",x"48"),
  1258 => (x"c3",x"c9",x"05",x"a8"),
  1259 => (x"a6",x"e4",x"c0",x"87"),
  1260 => (x"7e",x"78",x"c0",x"48"),
  1261 => (x"fb",x"c0",x"48",x"74"),
  1262 => (x"a6",x"ec",x"c0",x"88"),
  1263 => (x"02",x"98",x"70",x"58"),
  1264 => (x"48",x"87",x"c8",x"c8"),
  1265 => (x"ec",x"c0",x"88",x"cb"),
  1266 => (x"98",x"70",x"58",x"a6"),
  1267 => (x"87",x"d0",x"c1",x"02"),
  1268 => (x"c0",x"88",x"c9",x"48"),
  1269 => (x"70",x"58",x"a6",x"ec"),
  1270 => (x"d6",x"c3",x"02",x"98"),
  1271 => (x"88",x"c4",x"48",x"87"),
  1272 => (x"58",x"a6",x"ec",x"c0"),
  1273 => (x"d0",x"02",x"98",x"70"),
  1274 => (x"88",x"c1",x"48",x"87"),
  1275 => (x"58",x"a6",x"ec",x"c0"),
  1276 => (x"c2",x"02",x"98",x"70"),
  1277 => (x"cc",x"c7",x"87",x"fd"),
  1278 => (x"48",x"a6",x"d8",x"87"),
  1279 => (x"e2",x"78",x"f0",x"c0"),
  1280 => (x"4c",x"70",x"87",x"df"),
  1281 => (x"02",x"ac",x"ec",x"c0"),
  1282 => (x"dc",x"87",x"c3",x"c0"),
  1283 => (x"ec",x"c0",x"5c",x"a6"),
  1284 => (x"87",x"cc",x"02",x"ac"),
  1285 => (x"70",x"87",x"ca",x"e2"),
  1286 => (x"ac",x"ec",x"c0",x"4c"),
  1287 => (x"87",x"f4",x"ff",x"05"),
  1288 => (x"02",x"ac",x"ec",x"c0"),
  1289 => (x"e1",x"87",x"c3",x"c0"),
  1290 => (x"66",x"d8",x"87",x"f7"),
  1291 => (x"49",x"66",x"d4",x"1e"),
  1292 => (x"49",x"66",x"d4",x"1e"),
  1293 => (x"da",x"df",x"c1",x"1e"),
  1294 => (x"49",x"66",x"d4",x"1e"),
  1295 => (x"c0",x"87",x"ce",x"f7"),
  1296 => (x"dc",x"1e",x"ca",x"1e"),
  1297 => (x"91",x"cb",x"49",x"66"),
  1298 => (x"81",x"66",x"d8",x"c1"),
  1299 => (x"c4",x"48",x"a6",x"d8"),
  1300 => (x"66",x"d8",x"78",x"a1"),
  1301 => (x"cc",x"e2",x"49",x"bf"),
  1302 => (x"c0",x"86",x"d8",x"87"),
  1303 => (x"c1",x"06",x"a8",x"b7"),
  1304 => (x"1e",x"c1",x"87",x"c4"),
  1305 => (x"66",x"c8",x"1e",x"de"),
  1306 => (x"f8",x"e1",x"49",x"bf"),
  1307 => (x"70",x"86",x"c8",x"87"),
  1308 => (x"08",x"c0",x"48",x"49"),
  1309 => (x"58",x"a6",x"dc",x"88"),
  1310 => (x"06",x"a8",x"b7",x"c0"),
  1311 => (x"d8",x"87",x"e7",x"c0"),
  1312 => (x"b7",x"dd",x"48",x"66"),
  1313 => (x"87",x"de",x"03",x"a8"),
  1314 => (x"d8",x"49",x"bf",x"6e"),
  1315 => (x"e0",x"c0",x"81",x"66"),
  1316 => (x"49",x"66",x"d8",x"51"),
  1317 => (x"bf",x"6e",x"81",x"c1"),
  1318 => (x"51",x"c1",x"c2",x"81"),
  1319 => (x"c2",x"49",x"66",x"d8"),
  1320 => (x"81",x"bf",x"6e",x"81"),
  1321 => (x"66",x"cc",x"51",x"c0"),
  1322 => (x"d0",x"80",x"c1",x"48"),
  1323 => (x"7e",x"c1",x"58",x"a6"),
  1324 => (x"e2",x"87",x"d8",x"c4"),
  1325 => (x"a6",x"dc",x"87",x"de"),
  1326 => (x"87",x"d8",x"e2",x"58"),
  1327 => (x"58",x"a6",x"ec",x"c0"),
  1328 => (x"05",x"a8",x"ec",x"c0"),
  1329 => (x"c0",x"87",x"ca",x"c0"),
  1330 => (x"d8",x"48",x"a6",x"e8"),
  1331 => (x"c4",x"c0",x"78",x"66"),
  1332 => (x"cc",x"df",x"ff",x"87"),
  1333 => (x"49",x"66",x"c4",x"87"),
  1334 => (x"c0",x"c1",x"91",x"cb"),
  1335 => (x"80",x"71",x"48",x"66"),
  1336 => (x"4a",x"6e",x"7e",x"70"),
  1337 => (x"49",x"6e",x"82",x"c8"),
  1338 => (x"66",x"d8",x"81",x"ca"),
  1339 => (x"66",x"e8",x"c0",x"51"),
  1340 => (x"d8",x"81",x"c1",x"49"),
  1341 => (x"48",x"c1",x"89",x"66"),
  1342 => (x"49",x"70",x"30",x"71"),
  1343 => (x"97",x"71",x"89",x"c1"),
  1344 => (x"d1",x"ef",x"c2",x"7a"),
  1345 => (x"66",x"d8",x"49",x"bf"),
  1346 => (x"4a",x"6a",x"97",x"29"),
  1347 => (x"c0",x"98",x"71",x"48"),
  1348 => (x"6e",x"58",x"a6",x"f0"),
  1349 => (x"69",x"81",x"c4",x"49"),
  1350 => (x"66",x"e0",x"c0",x"4d"),
  1351 => (x"a8",x"66",x"dc",x"48"),
  1352 => (x"87",x"c8",x"c0",x"02"),
  1353 => (x"c0",x"48",x"a6",x"d8"),
  1354 => (x"87",x"c5",x"c0",x"78"),
  1355 => (x"c1",x"48",x"a6",x"d8"),
  1356 => (x"1e",x"66",x"d8",x"78"),
  1357 => (x"75",x"1e",x"e0",x"c0"),
  1358 => (x"e8",x"de",x"ff",x"49"),
  1359 => (x"70",x"86",x"c8",x"87"),
  1360 => (x"ac",x"b7",x"c0",x"4c"),
  1361 => (x"87",x"d4",x"c1",x"06"),
  1362 => (x"e0",x"c0",x"85",x"74"),
  1363 => (x"75",x"89",x"74",x"49"),
  1364 => (x"d6",x"d9",x"c1",x"4b"),
  1365 => (x"ed",x"fe",x"71",x"4a"),
  1366 => (x"85",x"c2",x"87",x"ce"),
  1367 => (x"48",x"66",x"e4",x"c0"),
  1368 => (x"e8",x"c0",x"80",x"c1"),
  1369 => (x"ec",x"c0",x"58",x"a6"),
  1370 => (x"81",x"c1",x"49",x"66"),
  1371 => (x"c0",x"02",x"a9",x"70"),
  1372 => (x"a6",x"d8",x"87",x"c8"),
  1373 => (x"c0",x"78",x"c0",x"48"),
  1374 => (x"a6",x"d8",x"87",x"c5"),
  1375 => (x"d8",x"78",x"c1",x"48"),
  1376 => (x"a4",x"c2",x"1e",x"66"),
  1377 => (x"48",x"e0",x"c0",x"49"),
  1378 => (x"49",x"70",x"88",x"71"),
  1379 => (x"ff",x"49",x"75",x"1e"),
  1380 => (x"c8",x"87",x"d2",x"dd"),
  1381 => (x"a8",x"b7",x"c0",x"86"),
  1382 => (x"87",x"c0",x"ff",x"01"),
  1383 => (x"02",x"66",x"e4",x"c0"),
  1384 => (x"6e",x"87",x"d1",x"c0"),
  1385 => (x"c0",x"81",x"c9",x"49"),
  1386 => (x"6e",x"51",x"66",x"e4"),
  1387 => (x"f9",x"c4",x"c1",x"48"),
  1388 => (x"87",x"cc",x"c0",x"78"),
  1389 => (x"81",x"c9",x"49",x"6e"),
  1390 => (x"48",x"6e",x"51",x"c2"),
  1391 => (x"78",x"ed",x"c5",x"c1"),
  1392 => (x"c6",x"c0",x"7e",x"c1"),
  1393 => (x"c8",x"dc",x"ff",x"87"),
  1394 => (x"6e",x"4c",x"70",x"87"),
  1395 => (x"87",x"f5",x"c0",x"02"),
  1396 => (x"c8",x"48",x"66",x"c4"),
  1397 => (x"c0",x"04",x"a8",x"66"),
  1398 => (x"66",x"c4",x"87",x"cb"),
  1399 => (x"c8",x"80",x"c1",x"48"),
  1400 => (x"e0",x"c0",x"58",x"a6"),
  1401 => (x"48",x"66",x"c8",x"87"),
  1402 => (x"a6",x"cc",x"88",x"c1"),
  1403 => (x"87",x"d5",x"c0",x"58"),
  1404 => (x"05",x"ac",x"c6",x"c1"),
  1405 => (x"cc",x"87",x"c8",x"c0"),
  1406 => (x"80",x"c1",x"48",x"66"),
  1407 => (x"ff",x"58",x"a6",x"d0"),
  1408 => (x"70",x"87",x"ce",x"db"),
  1409 => (x"48",x"66",x"d0",x"4c"),
  1410 => (x"a6",x"d4",x"80",x"c1"),
  1411 => (x"02",x"9c",x"74",x"58"),
  1412 => (x"c4",x"87",x"cb",x"c0"),
  1413 => (x"c8",x"c1",x"48",x"66"),
  1414 => (x"f3",x"04",x"a8",x"66"),
  1415 => (x"da",x"ff",x"87",x"d1"),
  1416 => (x"66",x"c4",x"87",x"e6"),
  1417 => (x"03",x"a8",x"c7",x"48"),
  1418 => (x"c2",x"87",x"e5",x"c0"),
  1419 => (x"c0",x"48",x"e4",x"eb"),
  1420 => (x"49",x"66",x"c4",x"78"),
  1421 => (x"c0",x"c1",x"91",x"cb"),
  1422 => (x"a1",x"c4",x"81",x"66"),
  1423 => (x"c0",x"4a",x"6a",x"4a"),
  1424 => (x"66",x"c4",x"79",x"52"),
  1425 => (x"c8",x"80",x"c1",x"48"),
  1426 => (x"a8",x"c7",x"58",x"a6"),
  1427 => (x"87",x"db",x"ff",x"04"),
  1428 => (x"e1",x"8e",x"d0",x"ff"),
  1429 => (x"20",x"3a",x"87",x"cd"),
  1430 => (x"1e",x"73",x"1e",x"00"),
  1431 => (x"02",x"9b",x"4b",x"71"),
  1432 => (x"eb",x"c2",x"87",x"c6"),
  1433 => (x"78",x"c0",x"48",x"e0"),
  1434 => (x"eb",x"c2",x"1e",x"c7"),
  1435 => (x"1e",x"49",x"bf",x"e0"),
  1436 => (x"1e",x"e7",x"dd",x"c1"),
  1437 => (x"bf",x"dc",x"eb",x"c2"),
  1438 => (x"87",x"c6",x"ef",x"49"),
  1439 => (x"eb",x"c2",x"86",x"cc"),
  1440 => (x"ea",x"49",x"bf",x"dc"),
  1441 => (x"9b",x"73",x"87",x"cb"),
  1442 => (x"c1",x"87",x"c8",x"02"),
  1443 => (x"c0",x"49",x"e7",x"dd"),
  1444 => (x"e0",x"87",x"d1",x"e7"),
  1445 => (x"73",x"1e",x"87",x"d1"),
  1446 => (x"c2",x"4b",x"c0",x"1e"),
  1447 => (x"c0",x"48",x"db",x"dc"),
  1448 => (x"ca",x"df",x"c1",x"50"),
  1449 => (x"fd",x"c0",x"49",x"bf"),
  1450 => (x"98",x"70",x"87",x"c6"),
  1451 => (x"c1",x"87",x"c4",x"05"),
  1452 => (x"73",x"4b",x"f9",x"da"),
  1453 => (x"ee",x"df",x"ff",x"48"),
  1454 => (x"4d",x"4f",x"52",x"87"),
  1455 => (x"61",x"6f",x"6c",x"20"),
  1456 => (x"67",x"6e",x"69",x"64"),
  1457 => (x"69",x"61",x"66",x"20"),
  1458 => (x"00",x"64",x"65",x"6c"),
  1459 => (x"87",x"e9",x"c7",x"1e"),
  1460 => (x"c4",x"fe",x"49",x"c1"),
  1461 => (x"e2",x"ef",x"fe",x"87"),
  1462 => (x"02",x"98",x"70",x"87"),
  1463 => (x"f8",x"fe",x"87",x"cd"),
  1464 => (x"98",x"70",x"87",x"df"),
  1465 => (x"c1",x"87",x"c4",x"02"),
  1466 => (x"c0",x"87",x"c2",x"4a"),
  1467 => (x"05",x"9a",x"72",x"4a"),
  1468 => (x"1e",x"c0",x"87",x"ce"),
  1469 => (x"49",x"e0",x"dc",x"c1"),
  1470 => (x"87",x"ed",x"f2",x"c0"),
  1471 => (x"87",x"fe",x"86",x"c4"),
  1472 => (x"87",x"c1",x"c1",x"c1"),
  1473 => (x"dc",x"c1",x"1e",x"c0"),
  1474 => (x"f2",x"c0",x"49",x"eb"),
  1475 => (x"1e",x"c0",x"87",x"db"),
  1476 => (x"70",x"87",x"c3",x"fe"),
  1477 => (x"d0",x"f2",x"c0",x"49"),
  1478 => (x"87",x"dc",x"c3",x"87"),
  1479 => (x"4f",x"26",x"8e",x"f8"),
  1480 => (x"66",x"20",x"44",x"53"),
  1481 => (x"65",x"6c",x"69",x"61"),
  1482 => (x"42",x"00",x"2e",x"64"),
  1483 => (x"69",x"74",x"6f",x"6f"),
  1484 => (x"2e",x"2e",x"67",x"6e"),
  1485 => (x"c0",x"1e",x"00",x"2e"),
  1486 => (x"c0",x"87",x"c5",x"e9"),
  1487 => (x"f6",x"87",x"e0",x"f5"),
  1488 => (x"1e",x"4f",x"26",x"87"),
  1489 => (x"48",x"e0",x"eb",x"c2"),
  1490 => (x"eb",x"c2",x"78",x"c0"),
  1491 => (x"78",x"c0",x"48",x"dc"),
  1492 => (x"e1",x"87",x"f9",x"fd"),
  1493 => (x"26",x"48",x"c0",x"87"),
  1494 => (x"45",x"20",x"80",x"4f"),
  1495 => (x"00",x"74",x"69",x"78"),
  1496 => (x"61",x"42",x"20",x"80"),
  1497 => (x"e9",x"00",x"6b",x"63"),
  1498 => (x"f5",x"00",x"00",x"10"),
  1499 => (x"00",x"00",x"00",x"2a"),
  1500 => (x"10",x"e9",x"00",x"00"),
  1501 => (x"2b",x"13",x"00",x"00"),
  1502 => (x"00",x"00",x"00",x"00"),
  1503 => (x"00",x"10",x"e9",x"00"),
  1504 => (x"00",x"2b",x"31",x"00"),
  1505 => (x"00",x"00",x"00",x"00"),
  1506 => (x"00",x"00",x"10",x"e9"),
  1507 => (x"00",x"00",x"2b",x"4f"),
  1508 => (x"e9",x"00",x"00",x"00"),
  1509 => (x"6d",x"00",x"00",x"10"),
  1510 => (x"00",x"00",x"00",x"2b"),
  1511 => (x"10",x"e9",x"00",x"00"),
  1512 => (x"2b",x"8b",x"00",x"00"),
  1513 => (x"00",x"00",x"00",x"00"),
  1514 => (x"00",x"10",x"e9",x"00"),
  1515 => (x"00",x"2b",x"a9",x"00"),
  1516 => (x"00",x"00",x"00",x"00"),
  1517 => (x"00",x"00",x"10",x"e9"),
  1518 => (x"00",x"00",x"00",x"00"),
  1519 => (x"7e",x"00",x"00",x"00"),
  1520 => (x"00",x"00",x"00",x"11"),
  1521 => (x"00",x"00",x"00",x"00"),
  1522 => (x"17",x"ce",x"00",x"00"),
  1523 => (x"45",x"4e",x"00",x"00"),
  1524 => (x"4f",x"45",x"47",x"4f"),
  1525 => (x"4f",x"52",x"20",x"20"),
  1526 => (x"6f",x"4c",x"00",x"4d"),
  1527 => (x"2a",x"20",x"64",x"61"),
  1528 => (x"fe",x"1e",x"00",x"2e"),
  1529 => (x"78",x"c0",x"48",x"f0"),
  1530 => (x"09",x"79",x"09",x"cd"),
  1531 => (x"1e",x"1e",x"4f",x"26"),
  1532 => (x"7e",x"bf",x"f0",x"fe"),
  1533 => (x"4f",x"26",x"26",x"48"),
  1534 => (x"48",x"f0",x"fe",x"1e"),
  1535 => (x"4f",x"26",x"78",x"c1"),
  1536 => (x"48",x"f0",x"fe",x"1e"),
  1537 => (x"4f",x"26",x"78",x"c0"),
  1538 => (x"c0",x"4a",x"71",x"1e"),
  1539 => (x"4f",x"26",x"52",x"52"),
  1540 => (x"5c",x"5b",x"5e",x"0e"),
  1541 => (x"86",x"f4",x"0e",x"5d"),
  1542 => (x"6d",x"97",x"4d",x"71"),
  1543 => (x"4c",x"a5",x"c1",x"7e"),
  1544 => (x"c8",x"48",x"6c",x"97"),
  1545 => (x"48",x"6e",x"58",x"a6"),
  1546 => (x"05",x"a8",x"66",x"c4"),
  1547 => (x"48",x"ff",x"87",x"c5"),
  1548 => (x"ff",x"87",x"e6",x"c0"),
  1549 => (x"a5",x"c2",x"87",x"ca"),
  1550 => (x"4b",x"6c",x"97",x"49"),
  1551 => (x"97",x"4b",x"a3",x"71"),
  1552 => (x"6c",x"97",x"4b",x"6b"),
  1553 => (x"c1",x"48",x"6e",x"7e"),
  1554 => (x"58",x"a6",x"c8",x"80"),
  1555 => (x"a6",x"cc",x"98",x"c7"),
  1556 => (x"7c",x"97",x"70",x"58"),
  1557 => (x"73",x"87",x"e1",x"fe"),
  1558 => (x"26",x"8e",x"f4",x"48"),
  1559 => (x"26",x"4c",x"26",x"4d"),
  1560 => (x"0e",x"4f",x"26",x"4b"),
  1561 => (x"0e",x"5c",x"5b",x"5e"),
  1562 => (x"4c",x"71",x"86",x"f4"),
  1563 => (x"c3",x"4a",x"66",x"d8"),
  1564 => (x"a4",x"c2",x"9a",x"ff"),
  1565 => (x"49",x"6c",x"97",x"4b"),
  1566 => (x"72",x"49",x"a1",x"73"),
  1567 => (x"7e",x"6c",x"97",x"51"),
  1568 => (x"80",x"c1",x"48",x"6e"),
  1569 => (x"c7",x"58",x"a6",x"c8"),
  1570 => (x"58",x"a6",x"cc",x"98"),
  1571 => (x"8e",x"f4",x"54",x"70"),
  1572 => (x"1e",x"87",x"ca",x"ff"),
  1573 => (x"87",x"e8",x"fd",x"1e"),
  1574 => (x"49",x"4a",x"bf",x"e0"),
  1575 => (x"99",x"c0",x"e0",x"c0"),
  1576 => (x"72",x"87",x"cb",x"02"),
  1577 => (x"c7",x"ef",x"c2",x"1e"),
  1578 => (x"87",x"f7",x"fe",x"49"),
  1579 => (x"fd",x"fc",x"86",x"c4"),
  1580 => (x"fd",x"7e",x"70",x"87"),
  1581 => (x"26",x"26",x"87",x"c2"),
  1582 => (x"ef",x"c2",x"1e",x"4f"),
  1583 => (x"c7",x"fd",x"49",x"c7"),
  1584 => (x"d3",x"e2",x"c1",x"87"),
  1585 => (x"87",x"da",x"fc",x"49"),
  1586 => (x"26",x"87",x"d5",x"c6"),
  1587 => (x"5b",x"5e",x"0e",x"4f"),
  1588 => (x"c2",x"0e",x"5d",x"5c"),
  1589 => (x"4a",x"bf",x"e6",x"ef"),
  1590 => (x"bf",x"e1",x"e4",x"c1"),
  1591 => (x"bc",x"72",x"4c",x"49"),
  1592 => (x"db",x"fc",x"4d",x"71"),
  1593 => (x"74",x"4b",x"c0",x"87"),
  1594 => (x"02",x"99",x"d0",x"49"),
  1595 => (x"49",x"75",x"87",x"d5"),
  1596 => (x"1e",x"71",x"99",x"d0"),
  1597 => (x"eb",x"c1",x"1e",x"c0"),
  1598 => (x"82",x"73",x"4a",x"ef"),
  1599 => (x"ca",x"c1",x"49",x"12"),
  1600 => (x"c1",x"86",x"c8",x"87"),
  1601 => (x"c8",x"83",x"2d",x"2c"),
  1602 => (x"da",x"ff",x"04",x"ab"),
  1603 => (x"87",x"e8",x"fb",x"87"),
  1604 => (x"48",x"e1",x"e4",x"c1"),
  1605 => (x"bf",x"e6",x"ef",x"c2"),
  1606 => (x"26",x"4d",x"26",x"78"),
  1607 => (x"26",x"4b",x"26",x"4c"),
  1608 => (x"00",x"00",x"00",x"4f"),
  1609 => (x"1e",x"73",x"1e",x"00"),
  1610 => (x"4a",x"c0",x"4b",x"71"),
  1611 => (x"49",x"ef",x"eb",x"c1"),
  1612 => (x"69",x"97",x"81",x"72"),
  1613 => (x"05",x"a9",x"73",x"49"),
  1614 => (x"48",x"c1",x"87",x"c4"),
  1615 => (x"82",x"c1",x"87",x"ca"),
  1616 => (x"04",x"aa",x"b7",x"c8"),
  1617 => (x"48",x"c0",x"87",x"e6"),
  1618 => (x"1e",x"87",x"d2",x"ff"),
  1619 => (x"4b",x"71",x"1e",x"73"),
  1620 => (x"87",x"d1",x"ff",x"49"),
  1621 => (x"c0",x"02",x"98",x"70"),
  1622 => (x"d0",x"ff",x"87",x"ec"),
  1623 => (x"78",x"e1",x"c8",x"48"),
  1624 => (x"c5",x"48",x"d4",x"ff"),
  1625 => (x"02",x"66",x"c8",x"78"),
  1626 => (x"e0",x"c3",x"87",x"c3"),
  1627 => (x"02",x"66",x"cc",x"78"),
  1628 => (x"d4",x"ff",x"87",x"c6"),
  1629 => (x"78",x"f0",x"c3",x"48"),
  1630 => (x"73",x"48",x"d4",x"ff"),
  1631 => (x"48",x"d0",x"ff",x"78"),
  1632 => (x"c0",x"78",x"e1",x"c8"),
  1633 => (x"d4",x"fe",x"78",x"e0"),
  1634 => (x"5b",x"5e",x"0e",x"87"),
  1635 => (x"4c",x"71",x"0e",x"5c"),
  1636 => (x"49",x"c7",x"ef",x"c2"),
  1637 => (x"70",x"87",x"f9",x"f9"),
  1638 => (x"aa",x"b7",x"c0",x"4a"),
  1639 => (x"87",x"e3",x"c2",x"04"),
  1640 => (x"05",x"aa",x"e0",x"c3"),
  1641 => (x"e9",x"c1",x"87",x"c9"),
  1642 => (x"78",x"c1",x"48",x"cc"),
  1643 => (x"c3",x"87",x"d4",x"c2"),
  1644 => (x"c9",x"05",x"aa",x"f0"),
  1645 => (x"c8",x"e9",x"c1",x"87"),
  1646 => (x"c1",x"78",x"c1",x"48"),
  1647 => (x"e9",x"c1",x"87",x"f5"),
  1648 => (x"c7",x"02",x"bf",x"cc"),
  1649 => (x"c2",x"4b",x"72",x"87"),
  1650 => (x"87",x"c2",x"b3",x"c0"),
  1651 => (x"9c",x"74",x"4b",x"72"),
  1652 => (x"c1",x"87",x"d1",x"05"),
  1653 => (x"1e",x"bf",x"c8",x"e9"),
  1654 => (x"bf",x"cc",x"e9",x"c1"),
  1655 => (x"fd",x"49",x"72",x"1e"),
  1656 => (x"86",x"c8",x"87",x"e9"),
  1657 => (x"bf",x"c8",x"e9",x"c1"),
  1658 => (x"87",x"e0",x"c0",x"02"),
  1659 => (x"b7",x"c4",x"49",x"73"),
  1660 => (x"ea",x"c1",x"91",x"29"),
  1661 => (x"4a",x"73",x"81",x"ef"),
  1662 => (x"92",x"c2",x"9a",x"cf"),
  1663 => (x"30",x"72",x"48",x"c1"),
  1664 => (x"ba",x"ff",x"4a",x"70"),
  1665 => (x"98",x"69",x"48",x"72"),
  1666 => (x"87",x"db",x"79",x"70"),
  1667 => (x"b7",x"c4",x"49",x"73"),
  1668 => (x"ea",x"c1",x"91",x"29"),
  1669 => (x"4a",x"73",x"81",x"ef"),
  1670 => (x"92",x"c2",x"9a",x"cf"),
  1671 => (x"30",x"72",x"48",x"c3"),
  1672 => (x"69",x"48",x"4a",x"70"),
  1673 => (x"c1",x"79",x"70",x"b0"),
  1674 => (x"c0",x"48",x"cc",x"e9"),
  1675 => (x"c8",x"e9",x"c1",x"78"),
  1676 => (x"c2",x"78",x"c0",x"48"),
  1677 => (x"f7",x"49",x"c7",x"ef"),
  1678 => (x"4a",x"70",x"87",x"d6"),
  1679 => (x"03",x"aa",x"b7",x"c0"),
  1680 => (x"c0",x"87",x"dd",x"fd"),
  1681 => (x"87",x"d3",x"fb",x"48"),
  1682 => (x"00",x"00",x"00",x"00"),
  1683 => (x"00",x"00",x"00",x"00"),
  1684 => (x"71",x"1e",x"73",x"1e"),
  1685 => (x"87",x"f5",x"f9",x"4b"),
  1686 => (x"ec",x"fc",x"49",x"73"),
  1687 => (x"87",x"fd",x"fa",x"87"),
  1688 => (x"72",x"4a",x"c0",x"1e"),
  1689 => (x"c1",x"91",x"c4",x"49"),
  1690 => (x"c0",x"81",x"ef",x"ea"),
  1691 => (x"d0",x"82",x"c1",x"79"),
  1692 => (x"ee",x"04",x"aa",x"b7"),
  1693 => (x"0e",x"4f",x"26",x"87"),
  1694 => (x"5d",x"5c",x"5b",x"5e"),
  1695 => (x"f5",x"4d",x"71",x"0e"),
  1696 => (x"4a",x"75",x"87",x"fe"),
  1697 => (x"92",x"2a",x"b7",x"c4"),
  1698 => (x"82",x"ef",x"ea",x"c1"),
  1699 => (x"9c",x"cf",x"4c",x"75"),
  1700 => (x"49",x"6a",x"94",x"c2"),
  1701 => (x"c3",x"2b",x"74",x"4b"),
  1702 => (x"74",x"48",x"c2",x"9b"),
  1703 => (x"ff",x"4c",x"70",x"30"),
  1704 => (x"71",x"48",x"74",x"bc"),
  1705 => (x"f5",x"7a",x"70",x"98"),
  1706 => (x"48",x"73",x"87",x"ce"),
  1707 => (x"00",x"87",x"ea",x"f9"),
  1708 => (x"00",x"00",x"00",x"00"),
  1709 => (x"00",x"00",x"00",x"00"),
  1710 => (x"00",x"00",x"00",x"00"),
  1711 => (x"00",x"00",x"00",x"00"),
  1712 => (x"00",x"00",x"00",x"00"),
  1713 => (x"00",x"00",x"00",x"00"),
  1714 => (x"00",x"00",x"00",x"00"),
  1715 => (x"00",x"00",x"00",x"00"),
  1716 => (x"00",x"00",x"00",x"00"),
  1717 => (x"00",x"00",x"00",x"00"),
  1718 => (x"00",x"00",x"00",x"00"),
  1719 => (x"00",x"00",x"00",x"00"),
  1720 => (x"00",x"00",x"00",x"00"),
  1721 => (x"00",x"00",x"00",x"00"),
  1722 => (x"00",x"00",x"00",x"00"),
  1723 => (x"16",x"00",x"00",x"00"),
  1724 => (x"2e",x"25",x"26",x"1e"),
  1725 => (x"1e",x"3e",x"3d",x"36"),
  1726 => (x"c8",x"48",x"d0",x"ff"),
  1727 => (x"48",x"71",x"78",x"e1"),
  1728 => (x"78",x"08",x"d4",x"ff"),
  1729 => (x"ff",x"1e",x"4f",x"26"),
  1730 => (x"e1",x"c8",x"48",x"d0"),
  1731 => (x"ff",x"48",x"71",x"78"),
  1732 => (x"c4",x"78",x"08",x"d4"),
  1733 => (x"d4",x"ff",x"48",x"66"),
  1734 => (x"4f",x"26",x"78",x"08"),
  1735 => (x"c4",x"4a",x"71",x"1e"),
  1736 => (x"72",x"1e",x"49",x"66"),
  1737 => (x"87",x"de",x"ff",x"49"),
  1738 => (x"c0",x"48",x"d0",x"ff"),
  1739 => (x"26",x"26",x"78",x"e0"),
  1740 => (x"4a",x"71",x"1e",x"4f"),
  1741 => (x"c1",x"1e",x"66",x"c4"),
  1742 => (x"ff",x"49",x"a2",x"e0"),
  1743 => (x"66",x"c8",x"87",x"c8"),
  1744 => (x"29",x"b7",x"c8",x"49"),
  1745 => (x"71",x"48",x"d4",x"ff"),
  1746 => (x"48",x"d0",x"ff",x"78"),
  1747 => (x"26",x"78",x"e0",x"c0"),
  1748 => (x"ff",x"1e",x"4f",x"26"),
  1749 => (x"ff",x"c3",x"4a",x"d4"),
  1750 => (x"48",x"d0",x"ff",x"7a"),
  1751 => (x"de",x"78",x"e1",x"c8"),
  1752 => (x"d1",x"ef",x"c2",x"7a"),
  1753 => (x"48",x"49",x"7a",x"bf"),
  1754 => (x"7a",x"70",x"28",x"c8"),
  1755 => (x"28",x"d0",x"48",x"71"),
  1756 => (x"48",x"71",x"7a",x"70"),
  1757 => (x"7a",x"70",x"28",x"d8"),
  1758 => (x"c0",x"48",x"d0",x"ff"),
  1759 => (x"4f",x"26",x"78",x"e0"),
  1760 => (x"5c",x"5b",x"5e",x"0e"),
  1761 => (x"4c",x"71",x"0e",x"5d"),
  1762 => (x"bf",x"d1",x"ef",x"c2"),
  1763 => (x"2b",x"74",x"4b",x"4d"),
  1764 => (x"c1",x"9b",x"66",x"d0"),
  1765 => (x"ab",x"66",x"d4",x"83"),
  1766 => (x"c0",x"87",x"c2",x"04"),
  1767 => (x"d0",x"4a",x"74",x"4b"),
  1768 => (x"31",x"72",x"49",x"66"),
  1769 => (x"99",x"75",x"b9",x"ff"),
  1770 => (x"30",x"72",x"48",x"73"),
  1771 => (x"71",x"48",x"4a",x"70"),
  1772 => (x"d5",x"ef",x"c2",x"b0"),
  1773 => (x"87",x"da",x"fe",x"58"),
  1774 => (x"4c",x"26",x"4d",x"26"),
  1775 => (x"4f",x"26",x"4b",x"26"),
  1776 => (x"48",x"d0",x"ff",x"1e"),
  1777 => (x"71",x"78",x"c9",x"c8"),
  1778 => (x"08",x"d4",x"ff",x"48"),
  1779 => (x"1e",x"4f",x"26",x"78"),
  1780 => (x"eb",x"49",x"4a",x"71"),
  1781 => (x"48",x"d0",x"ff",x"87"),
  1782 => (x"4f",x"26",x"78",x"c8"),
  1783 => (x"71",x"1e",x"73",x"1e"),
  1784 => (x"e1",x"ef",x"c2",x"4b"),
  1785 => (x"87",x"c3",x"02",x"bf"),
  1786 => (x"ff",x"87",x"eb",x"c2"),
  1787 => (x"c9",x"c8",x"48",x"d0"),
  1788 => (x"c0",x"49",x"73",x"78"),
  1789 => (x"d4",x"ff",x"b1",x"e0"),
  1790 => (x"c2",x"78",x"71",x"48"),
  1791 => (x"c0",x"48",x"d5",x"ef"),
  1792 => (x"02",x"66",x"c8",x"78"),
  1793 => (x"ff",x"c3",x"87",x"c5"),
  1794 => (x"c0",x"87",x"c2",x"49"),
  1795 => (x"dd",x"ef",x"c2",x"49"),
  1796 => (x"02",x"66",x"cc",x"59"),
  1797 => (x"d5",x"c5",x"87",x"c6"),
  1798 => (x"87",x"c4",x"4a",x"d5"),
  1799 => (x"4a",x"ff",x"ff",x"cf"),
  1800 => (x"5a",x"e1",x"ef",x"c2"),
  1801 => (x"48",x"e1",x"ef",x"c2"),
  1802 => (x"87",x"c4",x"78",x"c1"),
  1803 => (x"4c",x"26",x"4d",x"26"),
  1804 => (x"4f",x"26",x"4b",x"26"),
  1805 => (x"5c",x"5b",x"5e",x"0e"),
  1806 => (x"4a",x"71",x"0e",x"5d"),
  1807 => (x"bf",x"dd",x"ef",x"c2"),
  1808 => (x"02",x"9a",x"72",x"4c"),
  1809 => (x"c8",x"49",x"87",x"cb"),
  1810 => (x"d2",x"ef",x"c1",x"91"),
  1811 => (x"c4",x"83",x"71",x"4b"),
  1812 => (x"d2",x"f3",x"c1",x"87"),
  1813 => (x"13",x"4d",x"c0",x"4b"),
  1814 => (x"c2",x"99",x"74",x"49"),
  1815 => (x"b9",x"bf",x"d9",x"ef"),
  1816 => (x"71",x"48",x"d4",x"ff"),
  1817 => (x"2c",x"b7",x"c1",x"78"),
  1818 => (x"ad",x"b7",x"c8",x"85"),
  1819 => (x"c2",x"87",x"e8",x"04"),
  1820 => (x"48",x"bf",x"d5",x"ef"),
  1821 => (x"ef",x"c2",x"80",x"c8"),
  1822 => (x"ef",x"fe",x"58",x"d9"),
  1823 => (x"1e",x"73",x"1e",x"87"),
  1824 => (x"4a",x"13",x"4b",x"71"),
  1825 => (x"87",x"cb",x"02",x"9a"),
  1826 => (x"e7",x"fe",x"49",x"72"),
  1827 => (x"9a",x"4a",x"13",x"87"),
  1828 => (x"fe",x"87",x"f5",x"05"),
  1829 => (x"c2",x"1e",x"87",x"da"),
  1830 => (x"49",x"bf",x"d5",x"ef"),
  1831 => (x"48",x"d5",x"ef",x"c2"),
  1832 => (x"c4",x"78",x"a1",x"c1"),
  1833 => (x"03",x"a9",x"b7",x"c0"),
  1834 => (x"d4",x"ff",x"87",x"db"),
  1835 => (x"d9",x"ef",x"c2",x"48"),
  1836 => (x"ef",x"c2",x"78",x"bf"),
  1837 => (x"c2",x"49",x"bf",x"d5"),
  1838 => (x"c1",x"48",x"d5",x"ef"),
  1839 => (x"c0",x"c4",x"78",x"a1"),
  1840 => (x"e5",x"04",x"a9",x"b7"),
  1841 => (x"48",x"d0",x"ff",x"87"),
  1842 => (x"ef",x"c2",x"78",x"c8"),
  1843 => (x"78",x"c0",x"48",x"e1"),
  1844 => (x"00",x"00",x"4f",x"26"),
  1845 => (x"00",x"00",x"00",x"00"),
  1846 => (x"00",x"00",x"00",x"00"),
  1847 => (x"00",x"5f",x"5f",x"00"),
  1848 => (x"03",x"00",x"00",x"00"),
  1849 => (x"03",x"03",x"00",x"03"),
  1850 => (x"7f",x"14",x"00",x"00"),
  1851 => (x"7f",x"7f",x"14",x"7f"),
  1852 => (x"24",x"00",x"00",x"14"),
  1853 => (x"3a",x"6b",x"6b",x"2e"),
  1854 => (x"6a",x"4c",x"00",x"12"),
  1855 => (x"56",x"6c",x"18",x"36"),
  1856 => (x"7e",x"30",x"00",x"32"),
  1857 => (x"3a",x"77",x"59",x"4f"),
  1858 => (x"00",x"00",x"40",x"68"),
  1859 => (x"00",x"03",x"07",x"04"),
  1860 => (x"00",x"00",x"00",x"00"),
  1861 => (x"41",x"63",x"3e",x"1c"),
  1862 => (x"00",x"00",x"00",x"00"),
  1863 => (x"1c",x"3e",x"63",x"41"),
  1864 => (x"2a",x"08",x"00",x"00"),
  1865 => (x"3e",x"1c",x"1c",x"3e"),
  1866 => (x"08",x"00",x"08",x"2a"),
  1867 => (x"08",x"3e",x"3e",x"08"),
  1868 => (x"00",x"00",x"00",x"08"),
  1869 => (x"00",x"60",x"e0",x"80"),
  1870 => (x"08",x"00",x"00",x"00"),
  1871 => (x"08",x"08",x"08",x"08"),
  1872 => (x"00",x"00",x"00",x"08"),
  1873 => (x"00",x"60",x"60",x"00"),
  1874 => (x"60",x"40",x"00",x"00"),
  1875 => (x"06",x"0c",x"18",x"30"),
  1876 => (x"3e",x"00",x"01",x"03"),
  1877 => (x"7f",x"4d",x"59",x"7f"),
  1878 => (x"04",x"00",x"00",x"3e"),
  1879 => (x"00",x"7f",x"7f",x"06"),
  1880 => (x"42",x"00",x"00",x"00"),
  1881 => (x"4f",x"59",x"71",x"63"),
  1882 => (x"22",x"00",x"00",x"46"),
  1883 => (x"7f",x"49",x"49",x"63"),
  1884 => (x"1c",x"18",x"00",x"36"),
  1885 => (x"7f",x"7f",x"13",x"16"),
  1886 => (x"27",x"00",x"00",x"10"),
  1887 => (x"7d",x"45",x"45",x"67"),
  1888 => (x"3c",x"00",x"00",x"39"),
  1889 => (x"79",x"49",x"4b",x"7e"),
  1890 => (x"01",x"00",x"00",x"30"),
  1891 => (x"0f",x"79",x"71",x"01"),
  1892 => (x"36",x"00",x"00",x"07"),
  1893 => (x"7f",x"49",x"49",x"7f"),
  1894 => (x"06",x"00",x"00",x"36"),
  1895 => (x"3f",x"69",x"49",x"4f"),
  1896 => (x"00",x"00",x"00",x"1e"),
  1897 => (x"00",x"66",x"66",x"00"),
  1898 => (x"00",x"00",x"00",x"00"),
  1899 => (x"00",x"66",x"e6",x"80"),
  1900 => (x"08",x"00",x"00",x"00"),
  1901 => (x"22",x"14",x"14",x"08"),
  1902 => (x"14",x"00",x"00",x"22"),
  1903 => (x"14",x"14",x"14",x"14"),
  1904 => (x"22",x"00",x"00",x"14"),
  1905 => (x"08",x"14",x"14",x"22"),
  1906 => (x"02",x"00",x"00",x"08"),
  1907 => (x"0f",x"59",x"51",x"03"),
  1908 => (x"7f",x"3e",x"00",x"06"),
  1909 => (x"1f",x"55",x"5d",x"41"),
  1910 => (x"7e",x"00",x"00",x"1e"),
  1911 => (x"7f",x"09",x"09",x"7f"),
  1912 => (x"7f",x"00",x"00",x"7e"),
  1913 => (x"7f",x"49",x"49",x"7f"),
  1914 => (x"1c",x"00",x"00",x"36"),
  1915 => (x"41",x"41",x"63",x"3e"),
  1916 => (x"7f",x"00",x"00",x"41"),
  1917 => (x"3e",x"63",x"41",x"7f"),
  1918 => (x"7f",x"00",x"00",x"1c"),
  1919 => (x"41",x"49",x"49",x"7f"),
  1920 => (x"7f",x"00",x"00",x"41"),
  1921 => (x"01",x"09",x"09",x"7f"),
  1922 => (x"3e",x"00",x"00",x"01"),
  1923 => (x"7b",x"49",x"41",x"7f"),
  1924 => (x"7f",x"00",x"00",x"7a"),
  1925 => (x"7f",x"08",x"08",x"7f"),
  1926 => (x"00",x"00",x"00",x"7f"),
  1927 => (x"41",x"7f",x"7f",x"41"),
  1928 => (x"20",x"00",x"00",x"00"),
  1929 => (x"7f",x"40",x"40",x"60"),
  1930 => (x"7f",x"7f",x"00",x"3f"),
  1931 => (x"63",x"36",x"1c",x"08"),
  1932 => (x"7f",x"00",x"00",x"41"),
  1933 => (x"40",x"40",x"40",x"7f"),
  1934 => (x"7f",x"7f",x"00",x"40"),
  1935 => (x"7f",x"06",x"0c",x"06"),
  1936 => (x"7f",x"7f",x"00",x"7f"),
  1937 => (x"7f",x"18",x"0c",x"06"),
  1938 => (x"3e",x"00",x"00",x"7f"),
  1939 => (x"7f",x"41",x"41",x"7f"),
  1940 => (x"7f",x"00",x"00",x"3e"),
  1941 => (x"0f",x"09",x"09",x"7f"),
  1942 => (x"7f",x"3e",x"00",x"06"),
  1943 => (x"7e",x"7f",x"61",x"41"),
  1944 => (x"7f",x"00",x"00",x"40"),
  1945 => (x"7f",x"19",x"09",x"7f"),
  1946 => (x"26",x"00",x"00",x"66"),
  1947 => (x"7b",x"59",x"4d",x"6f"),
  1948 => (x"01",x"00",x"00",x"32"),
  1949 => (x"01",x"7f",x"7f",x"01"),
  1950 => (x"3f",x"00",x"00",x"01"),
  1951 => (x"7f",x"40",x"40",x"7f"),
  1952 => (x"0f",x"00",x"00",x"3f"),
  1953 => (x"3f",x"70",x"70",x"3f"),
  1954 => (x"7f",x"7f",x"00",x"0f"),
  1955 => (x"7f",x"30",x"18",x"30"),
  1956 => (x"63",x"41",x"00",x"7f"),
  1957 => (x"36",x"1c",x"1c",x"36"),
  1958 => (x"03",x"01",x"41",x"63"),
  1959 => (x"06",x"7c",x"7c",x"06"),
  1960 => (x"71",x"61",x"01",x"03"),
  1961 => (x"43",x"47",x"4d",x"59"),
  1962 => (x"00",x"00",x"00",x"41"),
  1963 => (x"41",x"41",x"7f",x"7f"),
  1964 => (x"03",x"01",x"00",x"00"),
  1965 => (x"30",x"18",x"0c",x"06"),
  1966 => (x"00",x"00",x"40",x"60"),
  1967 => (x"7f",x"7f",x"41",x"41"),
  1968 => (x"0c",x"08",x"00",x"00"),
  1969 => (x"0c",x"06",x"03",x"06"),
  1970 => (x"80",x"80",x"00",x"08"),
  1971 => (x"80",x"80",x"80",x"80"),
  1972 => (x"00",x"00",x"00",x"80"),
  1973 => (x"04",x"07",x"03",x"00"),
  1974 => (x"20",x"00",x"00",x"00"),
  1975 => (x"7c",x"54",x"54",x"74"),
  1976 => (x"7f",x"00",x"00",x"78"),
  1977 => (x"7c",x"44",x"44",x"7f"),
  1978 => (x"38",x"00",x"00",x"38"),
  1979 => (x"44",x"44",x"44",x"7c"),
  1980 => (x"38",x"00",x"00",x"00"),
  1981 => (x"7f",x"44",x"44",x"7c"),
  1982 => (x"38",x"00",x"00",x"7f"),
  1983 => (x"5c",x"54",x"54",x"7c"),
  1984 => (x"04",x"00",x"00",x"18"),
  1985 => (x"05",x"05",x"7f",x"7e"),
  1986 => (x"18",x"00",x"00",x"00"),
  1987 => (x"fc",x"a4",x"a4",x"bc"),
  1988 => (x"7f",x"00",x"00",x"7c"),
  1989 => (x"7c",x"04",x"04",x"7f"),
  1990 => (x"00",x"00",x"00",x"78"),
  1991 => (x"40",x"7d",x"3d",x"00"),
  1992 => (x"80",x"00",x"00",x"00"),
  1993 => (x"7d",x"fd",x"80",x"80"),
  1994 => (x"7f",x"00",x"00",x"00"),
  1995 => (x"6c",x"38",x"10",x"7f"),
  1996 => (x"00",x"00",x"00",x"44"),
  1997 => (x"40",x"7f",x"3f",x"00"),
  1998 => (x"7c",x"7c",x"00",x"00"),
  1999 => (x"7c",x"0c",x"18",x"0c"),
  2000 => (x"7c",x"00",x"00",x"78"),
  2001 => (x"7c",x"04",x"04",x"7c"),
  2002 => (x"38",x"00",x"00",x"78"),
  2003 => (x"7c",x"44",x"44",x"7c"),
  2004 => (x"fc",x"00",x"00",x"38"),
  2005 => (x"3c",x"24",x"24",x"fc"),
  2006 => (x"18",x"00",x"00",x"18"),
  2007 => (x"fc",x"24",x"24",x"3c"),
  2008 => (x"7c",x"00",x"00",x"fc"),
  2009 => (x"0c",x"04",x"04",x"7c"),
  2010 => (x"48",x"00",x"00",x"08"),
  2011 => (x"74",x"54",x"54",x"5c"),
  2012 => (x"04",x"00",x"00",x"20"),
  2013 => (x"44",x"44",x"7f",x"3f"),
  2014 => (x"3c",x"00",x"00",x"00"),
  2015 => (x"7c",x"40",x"40",x"7c"),
  2016 => (x"1c",x"00",x"00",x"7c"),
  2017 => (x"3c",x"60",x"60",x"3c"),
  2018 => (x"7c",x"3c",x"00",x"1c"),
  2019 => (x"7c",x"60",x"30",x"60"),
  2020 => (x"6c",x"44",x"00",x"3c"),
  2021 => (x"6c",x"38",x"10",x"38"),
  2022 => (x"1c",x"00",x"00",x"44"),
  2023 => (x"3c",x"60",x"e0",x"bc"),
  2024 => (x"44",x"00",x"00",x"1c"),
  2025 => (x"4c",x"5c",x"74",x"64"),
  2026 => (x"08",x"00",x"00",x"44"),
  2027 => (x"41",x"77",x"3e",x"08"),
  2028 => (x"00",x"00",x"00",x"41"),
  2029 => (x"00",x"7f",x"7f",x"00"),
  2030 => (x"41",x"00",x"00",x"00"),
  2031 => (x"08",x"3e",x"77",x"41"),
  2032 => (x"01",x"02",x"00",x"08"),
  2033 => (x"02",x"02",x"03",x"01"),
  2034 => (x"7f",x"7f",x"00",x"01"),
  2035 => (x"7f",x"7f",x"7f",x"7f"),
  2036 => (x"08",x"08",x"00",x"7f"),
  2037 => (x"3e",x"3e",x"1c",x"1c"),
  2038 => (x"7f",x"7f",x"7f",x"7f"),
  2039 => (x"1c",x"1c",x"3e",x"3e"),
  2040 => (x"10",x"00",x"08",x"08"),
  2041 => (x"18",x"7c",x"7c",x"18"),
  2042 => (x"10",x"00",x"00",x"10"),
  2043 => (x"30",x"7c",x"7c",x"30"),
  2044 => (x"30",x"10",x"00",x"10"),
  2045 => (x"1e",x"78",x"60",x"60"),
  2046 => (x"66",x"42",x"00",x"06"),
  2047 => (x"66",x"3c",x"18",x"3c"),
  2048 => (x"38",x"78",x"00",x"42"),
  2049 => (x"6c",x"c6",x"c2",x"6a"),
  2050 => (x"00",x"60",x"00",x"38"),
  2051 => (x"00",x"00",x"60",x"00"),
  2052 => (x"5e",x"0e",x"00",x"60"),
  2053 => (x"0e",x"5d",x"5c",x"5b"),
  2054 => (x"c2",x"4c",x"71",x"1e"),
  2055 => (x"4d",x"bf",x"f2",x"ef"),
  2056 => (x"1e",x"c0",x"4b",x"c0"),
  2057 => (x"c7",x"02",x"ab",x"74"),
  2058 => (x"48",x"a6",x"c4",x"87"),
  2059 => (x"87",x"c5",x"78",x"c0"),
  2060 => (x"c1",x"48",x"a6",x"c4"),
  2061 => (x"1e",x"66",x"c4",x"78"),
  2062 => (x"df",x"ee",x"49",x"73"),
  2063 => (x"c0",x"86",x"c8",x"87"),
  2064 => (x"ef",x"ef",x"49",x"e0"),
  2065 => (x"4a",x"a5",x"c4",x"87"),
  2066 => (x"f0",x"f0",x"49",x"6a"),
  2067 => (x"87",x"c6",x"f1",x"87"),
  2068 => (x"83",x"c1",x"85",x"cb"),
  2069 => (x"04",x"ab",x"b7",x"c8"),
  2070 => (x"26",x"87",x"c7",x"ff"),
  2071 => (x"4c",x"26",x"4d",x"26"),
  2072 => (x"4f",x"26",x"4b",x"26"),
  2073 => (x"c2",x"4a",x"71",x"1e"),
  2074 => (x"c2",x"5a",x"f6",x"ef"),
  2075 => (x"c7",x"48",x"f6",x"ef"),
  2076 => (x"dd",x"fe",x"49",x"78"),
  2077 => (x"1e",x"4f",x"26",x"87"),
  2078 => (x"4a",x"71",x"1e",x"73"),
  2079 => (x"03",x"aa",x"b7",x"c0"),
  2080 => (x"cf",x"c2",x"87",x"d3"),
  2081 => (x"c4",x"05",x"bf",x"fe"),
  2082 => (x"c2",x"4b",x"c1",x"87"),
  2083 => (x"c2",x"4b",x"c0",x"87"),
  2084 => (x"c4",x"5b",x"c2",x"d0"),
  2085 => (x"c2",x"d0",x"c2",x"87"),
  2086 => (x"fe",x"cf",x"c2",x"5a"),
  2087 => (x"9a",x"c1",x"4a",x"bf"),
  2088 => (x"49",x"a2",x"c0",x"c1"),
  2089 => (x"fc",x"87",x"e8",x"ec"),
  2090 => (x"fe",x"cf",x"c2",x"48"),
  2091 => (x"ef",x"fe",x"78",x"bf"),
  2092 => (x"4a",x"71",x"1e",x"87"),
  2093 => (x"72",x"1e",x"66",x"c4"),
  2094 => (x"87",x"f5",x"e9",x"49"),
  2095 => (x"1e",x"4f",x"26",x"26"),
  2096 => (x"bf",x"fe",x"cf",x"c2"),
  2097 => (x"87",x"c8",x"e6",x"49"),
  2098 => (x"48",x"ea",x"ef",x"c2"),
  2099 => (x"c2",x"78",x"bf",x"e8"),
  2100 => (x"ec",x"48",x"e6",x"ef"),
  2101 => (x"ef",x"c2",x"78",x"bf"),
  2102 => (x"49",x"4a",x"bf",x"ea"),
  2103 => (x"ca",x"99",x"ff",x"cf"),
  2104 => (x"48",x"72",x"2a",x"b7"),
  2105 => (x"ef",x"c2",x"b0",x"71"),
  2106 => (x"4f",x"26",x"58",x"f2"),
  2107 => (x"5c",x"5b",x"5e",x"0e"),
  2108 => (x"4b",x"71",x"0e",x"5d"),
  2109 => (x"c2",x"87",x"c8",x"ff"),
  2110 => (x"c0",x"48",x"e5",x"ef"),
  2111 => (x"e5",x"49",x"73",x"50"),
  2112 => (x"49",x"70",x"87",x"f5"),
  2113 => (x"cb",x"9c",x"c2",x"4c"),
  2114 => (x"f9",x"cb",x"49",x"ee"),
  2115 => (x"4d",x"49",x"70",x"87"),
  2116 => (x"97",x"e5",x"ef",x"c2"),
  2117 => (x"e2",x"c1",x"05",x"bf"),
  2118 => (x"49",x"66",x"d0",x"87"),
  2119 => (x"bf",x"ee",x"ef",x"c2"),
  2120 => (x"87",x"d6",x"05",x"99"),
  2121 => (x"c2",x"49",x"66",x"d4"),
  2122 => (x"99",x"bf",x"e6",x"ef"),
  2123 => (x"73",x"87",x"cb",x"05"),
  2124 => (x"87",x"c3",x"e5",x"49"),
  2125 => (x"c1",x"02",x"98",x"70"),
  2126 => (x"4c",x"c1",x"87",x"c1"),
  2127 => (x"75",x"87",x"c0",x"fe"),
  2128 => (x"87",x"ce",x"cb",x"49"),
  2129 => (x"c6",x"02",x"98",x"70"),
  2130 => (x"e5",x"ef",x"c2",x"87"),
  2131 => (x"c2",x"50",x"c1",x"48"),
  2132 => (x"bf",x"97",x"e5",x"ef"),
  2133 => (x"87",x"e3",x"c0",x"05"),
  2134 => (x"bf",x"ee",x"ef",x"c2"),
  2135 => (x"99",x"66",x"d0",x"49"),
  2136 => (x"87",x"d6",x"ff",x"05"),
  2137 => (x"bf",x"e6",x"ef",x"c2"),
  2138 => (x"99",x"66",x"d4",x"49"),
  2139 => (x"87",x"ca",x"ff",x"05"),
  2140 => (x"c2",x"e4",x"49",x"73"),
  2141 => (x"05",x"98",x"70",x"87"),
  2142 => (x"74",x"87",x"ff",x"fe"),
  2143 => (x"87",x"dc",x"fb",x"48"),
  2144 => (x"5c",x"5b",x"5e",x"0e"),
  2145 => (x"86",x"f4",x"0e",x"5d"),
  2146 => (x"ec",x"4c",x"4d",x"c0"),
  2147 => (x"a6",x"c4",x"7e",x"bf"),
  2148 => (x"f2",x"ef",x"c2",x"48"),
  2149 => (x"1e",x"c1",x"78",x"bf"),
  2150 => (x"49",x"c7",x"1e",x"c0"),
  2151 => (x"c8",x"87",x"cd",x"fd"),
  2152 => (x"02",x"98",x"70",x"86"),
  2153 => (x"49",x"ff",x"87",x"cd"),
  2154 => (x"c1",x"87",x"cc",x"fb"),
  2155 => (x"c6",x"e3",x"49",x"da"),
  2156 => (x"c2",x"4d",x"c1",x"87"),
  2157 => (x"bf",x"97",x"e5",x"ef"),
  2158 => (x"d5",x"87",x"c3",x"02"),
  2159 => (x"ef",x"c2",x"87",x"de"),
  2160 => (x"c2",x"4b",x"bf",x"ea"),
  2161 => (x"05",x"bf",x"fe",x"cf"),
  2162 => (x"c4",x"87",x"da",x"c1"),
  2163 => (x"c0",x"c2",x"48",x"a6"),
  2164 => (x"c2",x"78",x"c0",x"c0"),
  2165 => (x"6e",x"7e",x"ee",x"dd"),
  2166 => (x"6e",x"49",x"bf",x"97"),
  2167 => (x"70",x"80",x"c1",x"48"),
  2168 => (x"d2",x"e2",x"71",x"7e"),
  2169 => (x"02",x"98",x"70",x"87"),
  2170 => (x"66",x"c4",x"87",x"c3"),
  2171 => (x"48",x"66",x"c4",x"b3"),
  2172 => (x"c8",x"28",x"b7",x"c1"),
  2173 => (x"98",x"70",x"58",x"a6"),
  2174 => (x"87",x"db",x"ff",x"05"),
  2175 => (x"e1",x"49",x"fd",x"c3"),
  2176 => (x"fa",x"c3",x"87",x"f5"),
  2177 => (x"87",x"ef",x"e1",x"49"),
  2178 => (x"ff",x"cf",x"49",x"73"),
  2179 => (x"c0",x"1e",x"71",x"99"),
  2180 => (x"87",x"dd",x"fa",x"49"),
  2181 => (x"b7",x"ca",x"49",x"73"),
  2182 => (x"c1",x"1e",x"71",x"29"),
  2183 => (x"87",x"d1",x"fa",x"49"),
  2184 => (x"ff",x"c5",x"86",x"c8"),
  2185 => (x"ee",x"ef",x"c2",x"87"),
  2186 => (x"02",x"9b",x"4b",x"bf"),
  2187 => (x"cf",x"c2",x"87",x"dd"),
  2188 => (x"c7",x"49",x"bf",x"fa"),
  2189 => (x"98",x"70",x"87",x"dc"),
  2190 => (x"c0",x"87",x"c4",x"05"),
  2191 => (x"c2",x"87",x"d2",x"4b"),
  2192 => (x"c1",x"c7",x"49",x"e0"),
  2193 => (x"fe",x"cf",x"c2",x"87"),
  2194 => (x"c2",x"87",x"c6",x"58"),
  2195 => (x"c0",x"48",x"fa",x"cf"),
  2196 => (x"c2",x"49",x"73",x"78"),
  2197 => (x"87",x"cd",x"05",x"99"),
  2198 => (x"e0",x"49",x"eb",x"c3"),
  2199 => (x"49",x"70",x"87",x"d9"),
  2200 => (x"c2",x"02",x"99",x"c2"),
  2201 => (x"73",x"4c",x"fb",x"87"),
  2202 => (x"05",x"99",x"c1",x"49"),
  2203 => (x"f4",x"c3",x"87",x"cd"),
  2204 => (x"87",x"c3",x"e0",x"49"),
  2205 => (x"99",x"c2",x"49",x"70"),
  2206 => (x"fa",x"87",x"c2",x"02"),
  2207 => (x"c8",x"49",x"73",x"4c"),
  2208 => (x"87",x"ce",x"05",x"99"),
  2209 => (x"ff",x"49",x"f5",x"c3"),
  2210 => (x"70",x"87",x"ec",x"df"),
  2211 => (x"02",x"99",x"c2",x"49"),
  2212 => (x"ef",x"c2",x"87",x"d5"),
  2213 => (x"ca",x"02",x"bf",x"f6"),
  2214 => (x"88",x"c1",x"48",x"87"),
  2215 => (x"58",x"fa",x"ef",x"c2"),
  2216 => (x"ff",x"87",x"c2",x"c0"),
  2217 => (x"73",x"4d",x"c1",x"4c"),
  2218 => (x"05",x"99",x"c4",x"49"),
  2219 => (x"f2",x"c3",x"87",x"ce"),
  2220 => (x"c2",x"df",x"ff",x"49"),
  2221 => (x"c2",x"49",x"70",x"87"),
  2222 => (x"87",x"dc",x"02",x"99"),
  2223 => (x"bf",x"f6",x"ef",x"c2"),
  2224 => (x"b7",x"c7",x"48",x"7e"),
  2225 => (x"cb",x"c0",x"03",x"a8"),
  2226 => (x"c1",x"48",x"6e",x"87"),
  2227 => (x"fa",x"ef",x"c2",x"80"),
  2228 => (x"87",x"c2",x"c0",x"58"),
  2229 => (x"4d",x"c1",x"4c",x"fe"),
  2230 => (x"ff",x"49",x"fd",x"c3"),
  2231 => (x"70",x"87",x"d8",x"de"),
  2232 => (x"02",x"99",x"c2",x"49"),
  2233 => (x"c2",x"87",x"d5",x"c0"),
  2234 => (x"02",x"bf",x"f6",x"ef"),
  2235 => (x"c2",x"87",x"c9",x"c0"),
  2236 => (x"c0",x"48",x"f6",x"ef"),
  2237 => (x"87",x"c2",x"c0",x"78"),
  2238 => (x"4d",x"c1",x"4c",x"fd"),
  2239 => (x"ff",x"49",x"fa",x"c3"),
  2240 => (x"70",x"87",x"f4",x"dd"),
  2241 => (x"02",x"99",x"c2",x"49"),
  2242 => (x"c2",x"87",x"d9",x"c0"),
  2243 => (x"48",x"bf",x"f6",x"ef"),
  2244 => (x"03",x"a8",x"b7",x"c7"),
  2245 => (x"c2",x"87",x"c9",x"c0"),
  2246 => (x"c7",x"48",x"f6",x"ef"),
  2247 => (x"87",x"c2",x"c0",x"78"),
  2248 => (x"4d",x"c1",x"4c",x"fc"),
  2249 => (x"03",x"ac",x"b7",x"c0"),
  2250 => (x"c4",x"87",x"d1",x"c0"),
  2251 => (x"d8",x"c1",x"4a",x"66"),
  2252 => (x"c0",x"02",x"6a",x"82"),
  2253 => (x"4b",x"6a",x"87",x"c6"),
  2254 => (x"0f",x"73",x"49",x"74"),
  2255 => (x"f0",x"c3",x"1e",x"c0"),
  2256 => (x"49",x"da",x"c1",x"1e"),
  2257 => (x"c8",x"87",x"e5",x"f6"),
  2258 => (x"02",x"98",x"70",x"86"),
  2259 => (x"c8",x"87",x"e2",x"c0"),
  2260 => (x"ef",x"c2",x"48",x"a6"),
  2261 => (x"c8",x"78",x"bf",x"f6"),
  2262 => (x"91",x"cb",x"49",x"66"),
  2263 => (x"71",x"48",x"66",x"c4"),
  2264 => (x"6e",x"7e",x"70",x"80"),
  2265 => (x"c8",x"c0",x"02",x"bf"),
  2266 => (x"4b",x"bf",x"6e",x"87"),
  2267 => (x"73",x"49",x"66",x"c8"),
  2268 => (x"02",x"9d",x"75",x"0f"),
  2269 => (x"c2",x"87",x"c8",x"c0"),
  2270 => (x"49",x"bf",x"f6",x"ef"),
  2271 => (x"c2",x"87",x"d3",x"f2"),
  2272 => (x"02",x"bf",x"c2",x"d0"),
  2273 => (x"49",x"87",x"dd",x"c0"),
  2274 => (x"70",x"87",x"c7",x"c2"),
  2275 => (x"d3",x"c0",x"02",x"98"),
  2276 => (x"f6",x"ef",x"c2",x"87"),
  2277 => (x"f9",x"f1",x"49",x"bf"),
  2278 => (x"f3",x"49",x"c0",x"87"),
  2279 => (x"d0",x"c2",x"87",x"d9"),
  2280 => (x"78",x"c0",x"48",x"c2"),
  2281 => (x"f3",x"f2",x"8e",x"f4"),
  2282 => (x"5b",x"5e",x"0e",x"87"),
  2283 => (x"1e",x"0e",x"5d",x"5c"),
  2284 => (x"ef",x"c2",x"4c",x"71"),
  2285 => (x"c1",x"49",x"bf",x"f2"),
  2286 => (x"c1",x"4d",x"a1",x"cd"),
  2287 => (x"7e",x"69",x"81",x"d1"),
  2288 => (x"cf",x"02",x"9c",x"74"),
  2289 => (x"4b",x"a5",x"c4",x"87"),
  2290 => (x"ef",x"c2",x"7b",x"74"),
  2291 => (x"f2",x"49",x"bf",x"f2"),
  2292 => (x"7b",x"6e",x"87",x"d2"),
  2293 => (x"c4",x"05",x"9c",x"74"),
  2294 => (x"c2",x"4b",x"c0",x"87"),
  2295 => (x"73",x"4b",x"c1",x"87"),
  2296 => (x"87",x"d3",x"f2",x"49"),
  2297 => (x"c7",x"02",x"66",x"d4"),
  2298 => (x"87",x"da",x"49",x"87"),
  2299 => (x"87",x"c2",x"4a",x"70"),
  2300 => (x"d0",x"c2",x"4a",x"c0"),
  2301 => (x"f1",x"26",x"5a",x"c6"),
  2302 => (x"00",x"00",x"87",x"e2"),
  2303 => (x"00",x"00",x"00",x"00"),
  2304 => (x"00",x"00",x"00",x"00"),
  2305 => (x"71",x"1e",x"00",x"00"),
  2306 => (x"bf",x"c8",x"ff",x"4a"),
  2307 => (x"48",x"a1",x"72",x"49"),
  2308 => (x"ff",x"1e",x"4f",x"26"),
  2309 => (x"fe",x"89",x"bf",x"c8"),
  2310 => (x"c0",x"c0",x"c0",x"c0"),
  2311 => (x"c4",x"01",x"a9",x"c0"),
  2312 => (x"c2",x"4a",x"c0",x"87"),
  2313 => (x"72",x"4a",x"c1",x"87"),
  2314 => (x"0e",x"4f",x"26",x"48"),
  2315 => (x"5d",x"5c",x"5b",x"5e"),
  2316 => (x"ff",x"4b",x"71",x"0e"),
  2317 => (x"66",x"d0",x"4c",x"d4"),
  2318 => (x"d6",x"78",x"c0",x"48"),
  2319 => (x"f6",x"da",x"ff",x"49"),
  2320 => (x"7c",x"ff",x"c3",x"87"),
  2321 => (x"ff",x"c3",x"49",x"6c"),
  2322 => (x"49",x"4d",x"71",x"99"),
  2323 => (x"c1",x"99",x"f0",x"c3"),
  2324 => (x"cb",x"05",x"a9",x"e0"),
  2325 => (x"7c",x"ff",x"c3",x"87"),
  2326 => (x"98",x"c3",x"48",x"6c"),
  2327 => (x"78",x"08",x"66",x"d0"),
  2328 => (x"6c",x"7c",x"ff",x"c3"),
  2329 => (x"31",x"c8",x"49",x"4a"),
  2330 => (x"6c",x"7c",x"ff",x"c3"),
  2331 => (x"72",x"b2",x"71",x"4a"),
  2332 => (x"c3",x"31",x"c8",x"49"),
  2333 => (x"4a",x"6c",x"7c",x"ff"),
  2334 => (x"49",x"72",x"b2",x"71"),
  2335 => (x"ff",x"c3",x"31",x"c8"),
  2336 => (x"71",x"4a",x"6c",x"7c"),
  2337 => (x"48",x"d0",x"ff",x"b2"),
  2338 => (x"73",x"78",x"e0",x"c0"),
  2339 => (x"87",x"c2",x"02",x"9b"),
  2340 => (x"48",x"75",x"7b",x"72"),
  2341 => (x"4c",x"26",x"4d",x"26"),
  2342 => (x"4f",x"26",x"4b",x"26"),
  2343 => (x"0e",x"4f",x"26",x"1e"),
  2344 => (x"0e",x"5c",x"5b",x"5e"),
  2345 => (x"1e",x"76",x"86",x"f8"),
  2346 => (x"fd",x"49",x"a6",x"c8"),
  2347 => (x"86",x"c4",x"87",x"fd"),
  2348 => (x"48",x"6e",x"4b",x"70"),
  2349 => (x"c2",x"01",x"a8",x"c0"),
  2350 => (x"4a",x"73",x"87",x"f0"),
  2351 => (x"c1",x"9a",x"f0",x"c3"),
  2352 => (x"c7",x"02",x"aa",x"d0"),
  2353 => (x"aa",x"e0",x"c1",x"87"),
  2354 => (x"87",x"de",x"c2",x"05"),
  2355 => (x"99",x"c8",x"49",x"73"),
  2356 => (x"ff",x"87",x"c3",x"02"),
  2357 => (x"4c",x"73",x"87",x"c6"),
  2358 => (x"ac",x"c2",x"9c",x"c3"),
  2359 => (x"87",x"c2",x"c1",x"05"),
  2360 => (x"c9",x"49",x"66",x"c4"),
  2361 => (x"c4",x"1e",x"71",x"31"),
  2362 => (x"92",x"d4",x"4a",x"66"),
  2363 => (x"49",x"fa",x"ef",x"c2"),
  2364 => (x"d2",x"fe",x"81",x"72"),
  2365 => (x"49",x"d8",x"87",x"f9"),
  2366 => (x"87",x"fb",x"d7",x"ff"),
  2367 => (x"c2",x"1e",x"c0",x"c8"),
  2368 => (x"fd",x"49",x"ea",x"de"),
  2369 => (x"ff",x"87",x"d4",x"ef"),
  2370 => (x"e0",x"c0",x"48",x"d0"),
  2371 => (x"ea",x"de",x"c2",x"78"),
  2372 => (x"4a",x"66",x"cc",x"1e"),
  2373 => (x"ef",x"c2",x"92",x"d4"),
  2374 => (x"81",x"72",x"49",x"fa"),
  2375 => (x"87",x"cc",x"d1",x"fe"),
  2376 => (x"ac",x"c1",x"86",x"cc"),
  2377 => (x"87",x"c2",x"c1",x"05"),
  2378 => (x"c9",x"49",x"66",x"c4"),
  2379 => (x"c4",x"1e",x"71",x"31"),
  2380 => (x"92",x"d4",x"4a",x"66"),
  2381 => (x"49",x"fa",x"ef",x"c2"),
  2382 => (x"d1",x"fe",x"81",x"72"),
  2383 => (x"de",x"c2",x"87",x"f1"),
  2384 => (x"66",x"c8",x"1e",x"ea"),
  2385 => (x"c2",x"92",x"d4",x"4a"),
  2386 => (x"72",x"49",x"fa",x"ef"),
  2387 => (x"d8",x"cf",x"fe",x"81"),
  2388 => (x"ff",x"49",x"d7",x"87"),
  2389 => (x"c8",x"87",x"e0",x"d6"),
  2390 => (x"de",x"c2",x"1e",x"c0"),
  2391 => (x"ed",x"fd",x"49",x"ea"),
  2392 => (x"86",x"cc",x"87",x"e3"),
  2393 => (x"c0",x"48",x"d0",x"ff"),
  2394 => (x"8e",x"f8",x"78",x"e0"),
  2395 => (x"0e",x"87",x"e7",x"fc"),
  2396 => (x"5d",x"5c",x"5b",x"5e"),
  2397 => (x"4d",x"71",x"1e",x"0e"),
  2398 => (x"d4",x"4c",x"d4",x"ff"),
  2399 => (x"c3",x"48",x"7e",x"66"),
  2400 => (x"c5",x"06",x"a8",x"b7"),
  2401 => (x"c1",x"48",x"c0",x"87"),
  2402 => (x"49",x"75",x"87",x"e2"),
  2403 => (x"87",x"f0",x"df",x"fe"),
  2404 => (x"66",x"c4",x"1e",x"75"),
  2405 => (x"c2",x"93",x"d4",x"4b"),
  2406 => (x"73",x"83",x"fa",x"ef"),
  2407 => (x"ec",x"ca",x"fe",x"49"),
  2408 => (x"6b",x"83",x"c8",x"87"),
  2409 => (x"48",x"d0",x"ff",x"4b"),
  2410 => (x"dd",x"78",x"e1",x"c8"),
  2411 => (x"c3",x"49",x"73",x"7c"),
  2412 => (x"7c",x"71",x"99",x"ff"),
  2413 => (x"b7",x"c8",x"49",x"73"),
  2414 => (x"99",x"ff",x"c3",x"29"),
  2415 => (x"49",x"73",x"7c",x"71"),
  2416 => (x"c3",x"29",x"b7",x"d0"),
  2417 => (x"7c",x"71",x"99",x"ff"),
  2418 => (x"b7",x"d8",x"49",x"73"),
  2419 => (x"c0",x"7c",x"71",x"29"),
  2420 => (x"7c",x"7c",x"7c",x"7c"),
  2421 => (x"7c",x"7c",x"7c",x"7c"),
  2422 => (x"7c",x"7c",x"7c",x"7c"),
  2423 => (x"c4",x"78",x"e0",x"c0"),
  2424 => (x"49",x"dc",x"1e",x"66"),
  2425 => (x"87",x"f4",x"d4",x"ff"),
  2426 => (x"48",x"73",x"86",x"c8"),
  2427 => (x"87",x"e4",x"fa",x"26"),
  2428 => (x"5c",x"5b",x"5e",x"0e"),
  2429 => (x"71",x"1e",x"0e",x"5d"),
  2430 => (x"4b",x"d4",x"ff",x"7e"),
  2431 => (x"f0",x"c2",x"1e",x"6e"),
  2432 => (x"c9",x"fe",x"49",x"ce"),
  2433 => (x"86",x"c4",x"87",x"c7"),
  2434 => (x"02",x"9d",x"4d",x"70"),
  2435 => (x"c2",x"87",x"c3",x"c3"),
  2436 => (x"4c",x"bf",x"d6",x"f0"),
  2437 => (x"dd",x"fe",x"49",x"6e"),
  2438 => (x"d0",x"ff",x"87",x"e6"),
  2439 => (x"78",x"c5",x"c8",x"48"),
  2440 => (x"c0",x"7b",x"d6",x"c1"),
  2441 => (x"c1",x"7b",x"15",x"4a"),
  2442 => (x"b7",x"e0",x"c0",x"82"),
  2443 => (x"87",x"f5",x"04",x"aa"),
  2444 => (x"c4",x"48",x"d0",x"ff"),
  2445 => (x"78",x"c5",x"c8",x"78"),
  2446 => (x"c1",x"7b",x"d3",x"c1"),
  2447 => (x"74",x"78",x"c4",x"7b"),
  2448 => (x"fc",x"c1",x"02",x"9c"),
  2449 => (x"ea",x"de",x"c2",x"87"),
  2450 => (x"4d",x"c0",x"c8",x"7e"),
  2451 => (x"ac",x"b7",x"c0",x"8c"),
  2452 => (x"c8",x"87",x"c6",x"03"),
  2453 => (x"c0",x"4d",x"a4",x"c0"),
  2454 => (x"db",x"eb",x"c2",x"4c"),
  2455 => (x"d0",x"49",x"bf",x"97"),
  2456 => (x"87",x"d2",x"02",x"99"),
  2457 => (x"f0",x"c2",x"1e",x"c0"),
  2458 => (x"ca",x"fe",x"49",x"ce"),
  2459 => (x"86",x"c4",x"87",x"fb"),
  2460 => (x"c0",x"4a",x"49",x"70"),
  2461 => (x"de",x"c2",x"87",x"ef"),
  2462 => (x"f0",x"c2",x"1e",x"ea"),
  2463 => (x"ca",x"fe",x"49",x"ce"),
  2464 => (x"86",x"c4",x"87",x"e7"),
  2465 => (x"ff",x"4a",x"49",x"70"),
  2466 => (x"c5",x"c8",x"48",x"d0"),
  2467 => (x"7b",x"d4",x"c1",x"78"),
  2468 => (x"7b",x"bf",x"97",x"6e"),
  2469 => (x"80",x"c1",x"48",x"6e"),
  2470 => (x"8d",x"c1",x"7e",x"70"),
  2471 => (x"87",x"f0",x"ff",x"05"),
  2472 => (x"c4",x"48",x"d0",x"ff"),
  2473 => (x"05",x"9a",x"72",x"78"),
  2474 => (x"48",x"c0",x"87",x"c5"),
  2475 => (x"c1",x"87",x"e5",x"c0"),
  2476 => (x"ce",x"f0",x"c2",x"1e"),
  2477 => (x"cf",x"c8",x"fe",x"49"),
  2478 => (x"74",x"86",x"c4",x"87"),
  2479 => (x"c4",x"fe",x"05",x"9c"),
  2480 => (x"48",x"d0",x"ff",x"87"),
  2481 => (x"c1",x"78",x"c5",x"c8"),
  2482 => (x"7b",x"c0",x"7b",x"d3"),
  2483 => (x"48",x"c1",x"78",x"c4"),
  2484 => (x"48",x"c0",x"87",x"c2"),
  2485 => (x"26",x"4d",x"26",x"26"),
  2486 => (x"26",x"4b",x"26",x"4c"),
  2487 => (x"5b",x"5e",x"0e",x"4f"),
  2488 => (x"4b",x"71",x"0e",x"5c"),
  2489 => (x"d8",x"02",x"66",x"cc"),
  2490 => (x"f0",x"c0",x"4c",x"87"),
  2491 => (x"87",x"d8",x"02",x"8c"),
  2492 => (x"8a",x"c1",x"4a",x"74"),
  2493 => (x"8a",x"87",x"d1",x"02"),
  2494 => (x"8a",x"87",x"cd",x"02"),
  2495 => (x"d7",x"87",x"c9",x"02"),
  2496 => (x"fb",x"49",x"73",x"87"),
  2497 => (x"87",x"d0",x"87",x"ea"),
  2498 => (x"49",x"c0",x"1e",x"74"),
  2499 => (x"74",x"87",x"e0",x"f9"),
  2500 => (x"f9",x"49",x"73",x"1e"),
  2501 => (x"86",x"c8",x"87",x"d9"),
  2502 => (x"00",x"87",x"fc",x"fe"),
  2503 => (x"ea",x"dd",x"c2",x"1e"),
  2504 => (x"b9",x"c1",x"49",x"bf"),
  2505 => (x"59",x"ee",x"dd",x"c2"),
  2506 => (x"c3",x"48",x"d4",x"ff"),
  2507 => (x"d0",x"ff",x"78",x"ff"),
  2508 => (x"78",x"e1",x"c8",x"48"),
  2509 => (x"c1",x"48",x"d4",x"ff"),
  2510 => (x"71",x"31",x"c4",x"78"),
  2511 => (x"48",x"d0",x"ff",x"78"),
  2512 => (x"26",x"78",x"e0",x"c0"),
  2513 => (x"dd",x"c2",x"1e",x"4f"),
  2514 => (x"f0",x"c2",x"1e",x"de"),
  2515 => (x"c3",x"fe",x"49",x"ce"),
  2516 => (x"86",x"c4",x"87",x"fb"),
  2517 => (x"c3",x"02",x"98",x"70"),
  2518 => (x"87",x"c0",x"ff",x"87"),
  2519 => (x"35",x"31",x"4f",x"26"),
  2520 => (x"20",x"5a",x"48",x"4b"),
  2521 => (x"46",x"43",x"20",x"20"),
  2522 => (x"00",x"00",x"00",x"47"),
  2523 => (x"9f",x"1a",x"00",x"00"),
  2524 => (x"14",x"11",x"12",x"58"),
  2525 => (x"23",x"1c",x"1b",x"1d"),
  2526 => (x"59",x"5a",x"a7",x"4a"),
  2527 => (x"f2",x"f5",x"94",x"91"),
  2528 => (x"f2",x"f5",x"f4",x"eb"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

